// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : AIE.Axi4Module.Axi4Full.Stream2Axi4WriteMasterInterfaceAddFifo
// Git hash  : 6d1480269f65659931465c8b65ad201e15ffd506



module AIE.Axi4Module.Axi4Full.Stream2Axi4WriteMasterInterfaceAddFifo (
  input               s_axis_valid,
  output              s_axis_ready,
  input      [31:0]   s_axis_payload,
  output              m_axi_awvalid,
  input               m_axi_awready,
  output     [31:0]   m_axi_awaddr,
  output     [3:0]    m_axi_awregion,
  output     [7:0]    m_axi_awlen,
  output     [2:0]    m_axi_awsize,
  output     [1:0]    m_axi_awburst,
  output     [3:0]    m_axi_awcache,
  output     [3:0]    m_axi_awqos,
  output     [2:0]    m_axi_awprot,
  output              m_axi_wvalid,
  input               m_axi_wready,
  output     [31:0]   m_axi_wdata,
  output     [3:0]    m_axi_wstrb,
  output              m_axi_wlast,
  input               m_axi_bvalid,
  output              m_axi_bready,
  input      [1:0]    m_axi_bresp,
  output              m_axi_arvalid,
  input               m_axi_arready,
  output     [31:0]   m_axi_araddr,
  output     [3:0]    m_axi_arregion,
  output     [7:0]    m_axi_arlen,
  output     [2:0]    m_axi_arsize,
  output     [1:0]    m_axi_arburst,
  output     [3:0]    m_axi_arcache,
  output     [3:0]    m_axi_arqos,
  output     [2:0]    m_axi_arprot,
  input               m_axi_rvalid,
  output              m_axi_rready,
  input      [31:0]   m_axi_rdata,
  input      [1:0]    m_axi_rresp,
  input               m_axi_rlast,
  input               aresetn,
  input               aclk
);
  wire                axi4Interconnection_s_axis_ready;
  wire                axi4Interconnection_m_axi_arvalid;
  wire       [31:0]   axi4Interconnection_m_axi_araddr;
  wire       [3:0]    axi4Interconnection_m_axi_arregion;
  wire       [7:0]    axi4Interconnection_m_axi_arlen;
  wire       [2:0]    axi4Interconnection_m_axi_arsize;
  wire       [1:0]    axi4Interconnection_m_axi_arburst;
  wire       [3:0]    axi4Interconnection_m_axi_arcache;
  wire       [3:0]    axi4Interconnection_m_axi_arqos;
  wire       [2:0]    axi4Interconnection_m_axi_arprot;
  wire                axi4Interconnection_m_axi_awvalid;
  wire       [31:0]   axi4Interconnection_m_axi_awaddr;
  wire       [3:0]    axi4Interconnection_m_axi_awregion;
  wire       [7:0]    axi4Interconnection_m_axi_awlen;
  wire       [2:0]    axi4Interconnection_m_axi_awsize;
  wire       [1:0]    axi4Interconnection_m_axi_awburst;
  wire       [3:0]    axi4Interconnection_m_axi_awcache;
  wire       [3:0]    axi4Interconnection_m_axi_awqos;
  wire       [2:0]    axi4Interconnection_m_axi_awprot;
  wire                axi4Interconnection_m_axi_wvalid;
  wire       [31:0]   axi4Interconnection_m_axi_wdata;
  wire       [3:0]    axi4Interconnection_m_axi_wstrb;
  wire                axi4Interconnection_m_axi_wlast;
  wire                axi4Interconnection_m_axi_rready;
  wire                axi4Interconnection_m_axi_bready;
  wire                fifoInstance_io_push_ready;
  wire                fifoInstance_io_pop_valid;
  wire       [31:0]   fifoInstance_io_pop_payload;
  wire       [8:0]    fifoInstance_io_occupancy;
  wire       [8:0]    fifoInstance_io_availability;

  AIE.Axi4Module.Axi4Full.Stream2Axi4WriteMasterInterface axi4Interconnection (
    .s_axis_valid      (fifoInstance_io_pop_valid           ), //i
    .s_axis_ready      (axi4Interconnection_s_axis_ready    ), //o
    .s_axis_payload    (fifoInstance_io_pop_payload         ), //i
    .m_axi_awvalid     (axi4Interconnection_m_axi_awvalid   ), //o
    .m_axi_awready     (m_axi_awready                       ), //i
    .m_axi_awaddr      (axi4Interconnection_m_axi_awaddr    ), //o
    .m_axi_awregion    (axi4Interconnection_m_axi_awregion  ), //o
    .m_axi_awlen       (axi4Interconnection_m_axi_awlen     ), //o
    .m_axi_awsize      (axi4Interconnection_m_axi_awsize    ), //o
    .m_axi_awburst     (axi4Interconnection_m_axi_awburst   ), //o
    .m_axi_awcache     (axi4Interconnection_m_axi_awcache   ), //o
    .m_axi_awqos       (axi4Interconnection_m_axi_awqos     ), //o
    .m_axi_awprot      (axi4Interconnection_m_axi_awprot    ), //o
    .m_axi_wvalid      (axi4Interconnection_m_axi_wvalid    ), //o
    .m_axi_wready      (m_axi_wready                        ), //i
    .m_axi_wdata       (axi4Interconnection_m_axi_wdata     ), //o
    .m_axi_wstrb       (axi4Interconnection_m_axi_wstrb     ), //o
    .m_axi_wlast       (axi4Interconnection_m_axi_wlast     ), //o
    .m_axi_bvalid      (m_axi_bvalid                        ), //i
    .m_axi_bready      (axi4Interconnection_m_axi_bready    ), //o
    .m_axi_bresp       (m_axi_bresp                         ), //i
    .m_axi_arvalid     (axi4Interconnection_m_axi_arvalid   ), //o
    .m_axi_arready     (m_axi_arready                       ), //i
    .m_axi_araddr      (axi4Interconnection_m_axi_araddr    ), //o
    .m_axi_arregion    (axi4Interconnection_m_axi_arregion  ), //o
    .m_axi_arlen       (axi4Interconnection_m_axi_arlen     ), //o
    .m_axi_arsize      (axi4Interconnection_m_axi_arsize    ), //o
    .m_axi_arburst     (axi4Interconnection_m_axi_arburst   ), //o
    .m_axi_arcache     (axi4Interconnection_m_axi_arcache   ), //o
    .m_axi_arqos       (axi4Interconnection_m_axi_arqos     ), //o
    .m_axi_arprot      (axi4Interconnection_m_axi_arprot    ), //o
    .m_axi_rvalid      (m_axi_rvalid                        ), //i
    .m_axi_rready      (axi4Interconnection_m_axi_rready    ), //o
    .m_axi_rdata       (m_axi_rdata                         ), //i
    .m_axi_rresp       (m_axi_rresp                         ), //i
    .m_axi_rlast       (m_axi_rlast                         ), //i
    .aresetn           (aresetn                             ), //i
    .aclk              (aclk                                )  //i
  );
  StreamFifo fifoInstance (
    .io_push_valid      (s_axis_valid                      ), //i
    .io_push_ready      (fifoInstance_io_push_ready        ), //o
    .io_push_payload    (s_axis_payload                    ), //i
    .io_pop_valid       (fifoInstance_io_pop_valid         ), //o
    .io_pop_ready       (axi4Interconnection_s_axis_ready  ), //i
    .io_pop_payload     (fifoInstance_io_pop_payload       ), //o
    .io_flush           (1'b0                              ), //i
    .io_occupancy       (fifoInstance_io_occupancy         ), //o
    .io_availability    (fifoInstance_io_availability      ), //o
    .aclk               (aclk                              ), //i
    .aresetn            (aresetn                           )  //i
  );
  assign s_axis_ready = fifoInstance_io_push_ready;
  assign m_axi_arvalid = axi4Interconnection_m_axi_arvalid;
  assign m_axi_araddr = axi4Interconnection_m_axi_araddr;
  assign m_axi_arregion = axi4Interconnection_m_axi_arregion;
  assign m_axi_arlen = axi4Interconnection_m_axi_arlen;
  assign m_axi_arsize = axi4Interconnection_m_axi_arsize;
  assign m_axi_arburst = axi4Interconnection_m_axi_arburst;
  assign m_axi_arcache = axi4Interconnection_m_axi_arcache;
  assign m_axi_arqos = axi4Interconnection_m_axi_arqos;
  assign m_axi_arprot = axi4Interconnection_m_axi_arprot;
  assign m_axi_awvalid = axi4Interconnection_m_axi_awvalid;
  assign m_axi_awaddr = axi4Interconnection_m_axi_awaddr;
  assign m_axi_awregion = axi4Interconnection_m_axi_awregion;
  assign m_axi_awlen = axi4Interconnection_m_axi_awlen;
  assign m_axi_awsize = axi4Interconnection_m_axi_awsize;
  assign m_axi_awburst = axi4Interconnection_m_axi_awburst;
  assign m_axi_awcache = axi4Interconnection_m_axi_awcache;
  assign m_axi_awqos = axi4Interconnection_m_axi_awqos;
  assign m_axi_awprot = axi4Interconnection_m_axi_awprot;
  assign m_axi_wvalid = axi4Interconnection_m_axi_wvalid;
  assign m_axi_wdata = axi4Interconnection_m_axi_wdata;
  assign m_axi_wstrb = axi4Interconnection_m_axi_wstrb;
  assign m_axi_wlast = axi4Interconnection_m_axi_wlast;
  assign m_axi_rready = axi4Interconnection_m_axi_rready;
  assign m_axi_bready = axi4Interconnection_m_axi_bready;

endmodule

module StreamFifo (
  input               io_push_valid,
  output              io_push_ready,
  input      [31:0]   io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [31:0]   io_pop_payload,
  input               io_flush,
  output     [8:0]    io_occupancy,
  output     [8:0]    io_availability,
  input               aclk,
  input               aresetn
);
  reg        [31:0]   _zz_logic_ram_port0;
  wire       [7:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [7:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [7:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [7:0]    logic_pushPtr_valueNext;
  reg        [7:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [7:0]    logic_popPtr_valueNext;
  reg        [7:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l933;
  wire       [7:0]    logic_ptrDif;
  reg [31:0] logic_ram [0:255];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {7'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {7'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  always @(posedge aclk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge aclk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= io_push_payload;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 8'hff);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 8'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 8'hff);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 8'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l933 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge aclk or posedge aresetn) begin
    if(aresetn) begin
      logic_pushPtr_value <= 8'h0;
      logic_popPtr_value <= 8'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l933) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module AIE.Axi4Module.Axi4Full.Stream2Axi4WriteMasterInterface (
  input               s_axis_valid,
  output reg          s_axis_ready,
  input      [31:0]   s_axis_payload,
  output              m_axi_awvalid,
  input               m_axi_awready,
  output reg [31:0]   m_axi_awaddr,
  output     [3:0]    m_axi_awregion,
  output     [7:0]    m_axi_awlen,
  output     [2:0]    m_axi_awsize,
  output     [1:0]    m_axi_awburst,
  output     [3:0]    m_axi_awcache,
  output     [3:0]    m_axi_awqos,
  output     [2:0]    m_axi_awprot,
  output reg          m_axi_wvalid,
  input               m_axi_wready,
  output reg [31:0]   m_axi_wdata,
  output     [3:0]    m_axi_wstrb,
  output              m_axi_wlast,
  input               m_axi_bvalid,
  output              m_axi_bready,
  input      [1:0]    m_axi_bresp,
  output              m_axi_arvalid,
  input               m_axi_arready,
  output     [31:0]   m_axi_araddr,
  output     [3:0]    m_axi_arregion,
  output     [7:0]    m_axi_arlen,
  output     [2:0]    m_axi_arsize,
  output     [1:0]    m_axi_arburst,
  output     [3:0]    m_axi_arcache,
  output     [3:0]    m_axi_arqos,
  output     [2:0]    m_axi_arprot,
  input               m_axi_rvalid,
  output              m_axi_rready,
  input      [31:0]   m_axi_rdata,
  input      [1:0]    m_axi_rresp,
  input               m_axi_rlast,
  input               aresetn,
  input               aclk
);
  wire       [8:0]    _zz__zz_m_axi_wdata_1;
  wire       [0:0]    _zz__zz_m_axi_wdata_1_1;
  wire       [8:0]    _zz__zz_when_Axi4WriteMaster_l55_1;
  wire       [0:0]    _zz__zz_when_Axi4WriteMaster_l55_1_1;
  wire       [7:0]    _zz__zz_5;
  wire       [1:0]    _zz_Axi4Incr_alignMask;
  wire       [11:0]   _zz_Axi4Incr_base;
  wire       [11:0]   _zz_Axi4Incr_base_1;
  wire       [11:0]   _zz_Axi4Incr_baseIncr;
  wire       [2:0]    _zz_Axi4Incr_wrapCase_1;
  wire       [2:0]    _zz_Axi4Incr_wrapCase_2;
  reg        [11:0]   _zz_Axi4Incr_result;
  wire       [10:0]   _zz_Axi4Incr_result_1;
  wire       [0:0]    _zz_Axi4Incr_result_2;
  wire       [9:0]    _zz_Axi4Incr_result_3;
  wire       [1:0]    _zz_Axi4Incr_result_4;
  wire       [8:0]    _zz_Axi4Incr_result_5;
  wire       [2:0]    _zz_Axi4Incr_result_6;
  wire       [7:0]    _zz_Axi4Incr_result_7;
  wire       [3:0]    _zz_Axi4Incr_result_8;
  wire       [6:0]    _zz_Axi4Incr_result_9;
  wire       [4:0]    _zz_Axi4Incr_result_10;
  wire       [5:0]    _zz_Axi4Incr_result_11;
  wire       [5:0]    _zz_Axi4Incr_result_12;
  reg        [31:0]   _zz_m_axi_wdata_3;
  wire       [7:0]    _zz_m_axi_wdata_4;
  reg                 _zz_m_axi_wdata;
  reg                 _zz_1;
  reg        [8:0]    _zz_m_axi_wdata_1;
  reg        [8:0]    _zz_m_axi_wdata_2;
  wire                _zz_when_Axi4WriteMaster_l92;
  wire                _zz_2;
  reg                 _zz_when_Axi4WriteMaster_l55;
  reg                 _zz_3;
  reg        [8:0]    _zz_when_Axi4WriteMaster_l55_1;
  reg        [8:0]    _zz_when_Axi4WriteMaster_l55_2;
  wire                _zz_when_Axi4WriteMaster_l55_3;
  wire                _zz_4;
  reg        [31:0]   axi4Interface_fifoDataBuffer_0;
  reg        [31:0]   axi4Interface_fifoDataBuffer_1;
  reg        [31:0]   axi4Interface_fifoDataBuffer_2;
  reg        [31:0]   axi4Interface_fifoDataBuffer_3;
  reg        [31:0]   axi4Interface_fifoDataBuffer_4;
  reg        [31:0]   axi4Interface_fifoDataBuffer_5;
  reg        [31:0]   axi4Interface_fifoDataBuffer_6;
  reg        [31:0]   axi4Interface_fifoDataBuffer_7;
  reg        [31:0]   axi4Interface_fifoDataBuffer_8;
  reg        [31:0]   axi4Interface_fifoDataBuffer_9;
  reg        [31:0]   axi4Interface_fifoDataBuffer_10;
  reg        [31:0]   axi4Interface_fifoDataBuffer_11;
  reg        [31:0]   axi4Interface_fifoDataBuffer_12;
  reg        [31:0]   axi4Interface_fifoDataBuffer_13;
  reg        [31:0]   axi4Interface_fifoDataBuffer_14;
  reg        [31:0]   axi4Interface_fifoDataBuffer_15;
  reg        [31:0]   axi4Interface_fifoDataBuffer_16;
  reg        [31:0]   axi4Interface_fifoDataBuffer_17;
  reg        [31:0]   axi4Interface_fifoDataBuffer_18;
  reg        [31:0]   axi4Interface_fifoDataBuffer_19;
  reg        [31:0]   axi4Interface_fifoDataBuffer_20;
  reg        [31:0]   axi4Interface_fifoDataBuffer_21;
  reg        [31:0]   axi4Interface_fifoDataBuffer_22;
  reg        [31:0]   axi4Interface_fifoDataBuffer_23;
  reg        [31:0]   axi4Interface_fifoDataBuffer_24;
  reg        [31:0]   axi4Interface_fifoDataBuffer_25;
  reg        [31:0]   axi4Interface_fifoDataBuffer_26;
  reg        [31:0]   axi4Interface_fifoDataBuffer_27;
  reg        [31:0]   axi4Interface_fifoDataBuffer_28;
  reg        [31:0]   axi4Interface_fifoDataBuffer_29;
  reg        [31:0]   axi4Interface_fifoDataBuffer_30;
  reg        [31:0]   axi4Interface_fifoDataBuffer_31;
  reg        [31:0]   axi4Interface_fifoDataBuffer_32;
  reg        [31:0]   axi4Interface_fifoDataBuffer_33;
  reg        [31:0]   axi4Interface_fifoDataBuffer_34;
  reg        [31:0]   axi4Interface_fifoDataBuffer_35;
  reg        [31:0]   axi4Interface_fifoDataBuffer_36;
  reg        [31:0]   axi4Interface_fifoDataBuffer_37;
  reg        [31:0]   axi4Interface_fifoDataBuffer_38;
  reg        [31:0]   axi4Interface_fifoDataBuffer_39;
  reg        [31:0]   axi4Interface_fifoDataBuffer_40;
  reg        [31:0]   axi4Interface_fifoDataBuffer_41;
  reg        [31:0]   axi4Interface_fifoDataBuffer_42;
  reg        [31:0]   axi4Interface_fifoDataBuffer_43;
  reg        [31:0]   axi4Interface_fifoDataBuffer_44;
  reg        [31:0]   axi4Interface_fifoDataBuffer_45;
  reg        [31:0]   axi4Interface_fifoDataBuffer_46;
  reg        [31:0]   axi4Interface_fifoDataBuffer_47;
  reg        [31:0]   axi4Interface_fifoDataBuffer_48;
  reg        [31:0]   axi4Interface_fifoDataBuffer_49;
  reg        [31:0]   axi4Interface_fifoDataBuffer_50;
  reg        [31:0]   axi4Interface_fifoDataBuffer_51;
  reg        [31:0]   axi4Interface_fifoDataBuffer_52;
  reg        [31:0]   axi4Interface_fifoDataBuffer_53;
  reg        [31:0]   axi4Interface_fifoDataBuffer_54;
  reg        [31:0]   axi4Interface_fifoDataBuffer_55;
  reg        [31:0]   axi4Interface_fifoDataBuffer_56;
  reg        [31:0]   axi4Interface_fifoDataBuffer_57;
  reg        [31:0]   axi4Interface_fifoDataBuffer_58;
  reg        [31:0]   axi4Interface_fifoDataBuffer_59;
  reg        [31:0]   axi4Interface_fifoDataBuffer_60;
  reg        [31:0]   axi4Interface_fifoDataBuffer_61;
  reg        [31:0]   axi4Interface_fifoDataBuffer_62;
  reg        [31:0]   axi4Interface_fifoDataBuffer_63;
  reg        [31:0]   axi4Interface_fifoDataBuffer_64;
  reg        [31:0]   axi4Interface_fifoDataBuffer_65;
  reg        [31:0]   axi4Interface_fifoDataBuffer_66;
  reg        [31:0]   axi4Interface_fifoDataBuffer_67;
  reg        [31:0]   axi4Interface_fifoDataBuffer_68;
  reg        [31:0]   axi4Interface_fifoDataBuffer_69;
  reg        [31:0]   axi4Interface_fifoDataBuffer_70;
  reg        [31:0]   axi4Interface_fifoDataBuffer_71;
  reg        [31:0]   axi4Interface_fifoDataBuffer_72;
  reg        [31:0]   axi4Interface_fifoDataBuffer_73;
  reg        [31:0]   axi4Interface_fifoDataBuffer_74;
  reg        [31:0]   axi4Interface_fifoDataBuffer_75;
  reg        [31:0]   axi4Interface_fifoDataBuffer_76;
  reg        [31:0]   axi4Interface_fifoDataBuffer_77;
  reg        [31:0]   axi4Interface_fifoDataBuffer_78;
  reg        [31:0]   axi4Interface_fifoDataBuffer_79;
  reg        [31:0]   axi4Interface_fifoDataBuffer_80;
  reg        [31:0]   axi4Interface_fifoDataBuffer_81;
  reg        [31:0]   axi4Interface_fifoDataBuffer_82;
  reg        [31:0]   axi4Interface_fifoDataBuffer_83;
  reg        [31:0]   axi4Interface_fifoDataBuffer_84;
  reg        [31:0]   axi4Interface_fifoDataBuffer_85;
  reg        [31:0]   axi4Interface_fifoDataBuffer_86;
  reg        [31:0]   axi4Interface_fifoDataBuffer_87;
  reg        [31:0]   axi4Interface_fifoDataBuffer_88;
  reg        [31:0]   axi4Interface_fifoDataBuffer_89;
  reg        [31:0]   axi4Interface_fifoDataBuffer_90;
  reg        [31:0]   axi4Interface_fifoDataBuffer_91;
  reg        [31:0]   axi4Interface_fifoDataBuffer_92;
  reg        [31:0]   axi4Interface_fifoDataBuffer_93;
  reg        [31:0]   axi4Interface_fifoDataBuffer_94;
  reg        [31:0]   axi4Interface_fifoDataBuffer_95;
  reg        [31:0]   axi4Interface_fifoDataBuffer_96;
  reg        [31:0]   axi4Interface_fifoDataBuffer_97;
  reg        [31:0]   axi4Interface_fifoDataBuffer_98;
  reg        [31:0]   axi4Interface_fifoDataBuffer_99;
  reg        [31:0]   axi4Interface_fifoDataBuffer_100;
  reg        [31:0]   axi4Interface_fifoDataBuffer_101;
  reg        [31:0]   axi4Interface_fifoDataBuffer_102;
  reg        [31:0]   axi4Interface_fifoDataBuffer_103;
  reg        [31:0]   axi4Interface_fifoDataBuffer_104;
  reg        [31:0]   axi4Interface_fifoDataBuffer_105;
  reg        [31:0]   axi4Interface_fifoDataBuffer_106;
  reg        [31:0]   axi4Interface_fifoDataBuffer_107;
  reg        [31:0]   axi4Interface_fifoDataBuffer_108;
  reg        [31:0]   axi4Interface_fifoDataBuffer_109;
  reg        [31:0]   axi4Interface_fifoDataBuffer_110;
  reg        [31:0]   axi4Interface_fifoDataBuffer_111;
  reg        [31:0]   axi4Interface_fifoDataBuffer_112;
  reg        [31:0]   axi4Interface_fifoDataBuffer_113;
  reg        [31:0]   axi4Interface_fifoDataBuffer_114;
  reg        [31:0]   axi4Interface_fifoDataBuffer_115;
  reg        [31:0]   axi4Interface_fifoDataBuffer_116;
  reg        [31:0]   axi4Interface_fifoDataBuffer_117;
  reg        [31:0]   axi4Interface_fifoDataBuffer_118;
  reg        [31:0]   axi4Interface_fifoDataBuffer_119;
  reg        [31:0]   axi4Interface_fifoDataBuffer_120;
  reg        [31:0]   axi4Interface_fifoDataBuffer_121;
  reg        [31:0]   axi4Interface_fifoDataBuffer_122;
  reg        [31:0]   axi4Interface_fifoDataBuffer_123;
  reg        [31:0]   axi4Interface_fifoDataBuffer_124;
  reg        [31:0]   axi4Interface_fifoDataBuffer_125;
  reg        [31:0]   axi4Interface_fifoDataBuffer_126;
  reg        [31:0]   axi4Interface_fifoDataBuffer_127;
  reg        [31:0]   axi4Interface_fifoDataBuffer_128;
  reg        [31:0]   axi4Interface_fifoDataBuffer_129;
  reg        [31:0]   axi4Interface_fifoDataBuffer_130;
  reg        [31:0]   axi4Interface_fifoDataBuffer_131;
  reg        [31:0]   axi4Interface_fifoDataBuffer_132;
  reg        [31:0]   axi4Interface_fifoDataBuffer_133;
  reg        [31:0]   axi4Interface_fifoDataBuffer_134;
  reg        [31:0]   axi4Interface_fifoDataBuffer_135;
  reg        [31:0]   axi4Interface_fifoDataBuffer_136;
  reg        [31:0]   axi4Interface_fifoDataBuffer_137;
  reg        [31:0]   axi4Interface_fifoDataBuffer_138;
  reg        [31:0]   axi4Interface_fifoDataBuffer_139;
  reg        [31:0]   axi4Interface_fifoDataBuffer_140;
  reg        [31:0]   axi4Interface_fifoDataBuffer_141;
  reg        [31:0]   axi4Interface_fifoDataBuffer_142;
  reg        [31:0]   axi4Interface_fifoDataBuffer_143;
  reg        [31:0]   axi4Interface_fifoDataBuffer_144;
  reg        [31:0]   axi4Interface_fifoDataBuffer_145;
  reg        [31:0]   axi4Interface_fifoDataBuffer_146;
  reg        [31:0]   axi4Interface_fifoDataBuffer_147;
  reg        [31:0]   axi4Interface_fifoDataBuffer_148;
  reg        [31:0]   axi4Interface_fifoDataBuffer_149;
  reg        [31:0]   axi4Interface_fifoDataBuffer_150;
  reg        [31:0]   axi4Interface_fifoDataBuffer_151;
  reg        [31:0]   axi4Interface_fifoDataBuffer_152;
  reg        [31:0]   axi4Interface_fifoDataBuffer_153;
  reg        [31:0]   axi4Interface_fifoDataBuffer_154;
  reg        [31:0]   axi4Interface_fifoDataBuffer_155;
  reg        [31:0]   axi4Interface_fifoDataBuffer_156;
  reg        [31:0]   axi4Interface_fifoDataBuffer_157;
  reg        [31:0]   axi4Interface_fifoDataBuffer_158;
  reg        [31:0]   axi4Interface_fifoDataBuffer_159;
  reg        [31:0]   axi4Interface_fifoDataBuffer_160;
  reg        [31:0]   axi4Interface_fifoDataBuffer_161;
  reg        [31:0]   axi4Interface_fifoDataBuffer_162;
  reg        [31:0]   axi4Interface_fifoDataBuffer_163;
  reg        [31:0]   axi4Interface_fifoDataBuffer_164;
  reg        [31:0]   axi4Interface_fifoDataBuffer_165;
  reg        [31:0]   axi4Interface_fifoDataBuffer_166;
  reg        [31:0]   axi4Interface_fifoDataBuffer_167;
  reg        [31:0]   axi4Interface_fifoDataBuffer_168;
  reg        [31:0]   axi4Interface_fifoDataBuffer_169;
  reg        [31:0]   axi4Interface_fifoDataBuffer_170;
  reg        [31:0]   axi4Interface_fifoDataBuffer_171;
  reg        [31:0]   axi4Interface_fifoDataBuffer_172;
  reg        [31:0]   axi4Interface_fifoDataBuffer_173;
  reg        [31:0]   axi4Interface_fifoDataBuffer_174;
  reg        [31:0]   axi4Interface_fifoDataBuffer_175;
  reg        [31:0]   axi4Interface_fifoDataBuffer_176;
  reg        [31:0]   axi4Interface_fifoDataBuffer_177;
  reg        [31:0]   axi4Interface_fifoDataBuffer_178;
  reg        [31:0]   axi4Interface_fifoDataBuffer_179;
  reg        [31:0]   axi4Interface_fifoDataBuffer_180;
  reg        [31:0]   axi4Interface_fifoDataBuffer_181;
  reg        [31:0]   axi4Interface_fifoDataBuffer_182;
  reg        [31:0]   axi4Interface_fifoDataBuffer_183;
  reg        [31:0]   axi4Interface_fifoDataBuffer_184;
  reg        [31:0]   axi4Interface_fifoDataBuffer_185;
  reg        [31:0]   axi4Interface_fifoDataBuffer_186;
  reg        [31:0]   axi4Interface_fifoDataBuffer_187;
  reg        [31:0]   axi4Interface_fifoDataBuffer_188;
  reg        [31:0]   axi4Interface_fifoDataBuffer_189;
  reg        [31:0]   axi4Interface_fifoDataBuffer_190;
  reg        [31:0]   axi4Interface_fifoDataBuffer_191;
  reg        [31:0]   axi4Interface_fifoDataBuffer_192;
  reg        [31:0]   axi4Interface_fifoDataBuffer_193;
  reg        [31:0]   axi4Interface_fifoDataBuffer_194;
  reg        [31:0]   axi4Interface_fifoDataBuffer_195;
  reg        [31:0]   axi4Interface_fifoDataBuffer_196;
  reg        [31:0]   axi4Interface_fifoDataBuffer_197;
  reg        [31:0]   axi4Interface_fifoDataBuffer_198;
  reg        [31:0]   axi4Interface_fifoDataBuffer_199;
  reg        [31:0]   axi4Interface_fifoDataBuffer_200;
  reg        [31:0]   axi4Interface_fifoDataBuffer_201;
  reg        [31:0]   axi4Interface_fifoDataBuffer_202;
  reg        [31:0]   axi4Interface_fifoDataBuffer_203;
  reg        [31:0]   axi4Interface_fifoDataBuffer_204;
  reg        [31:0]   axi4Interface_fifoDataBuffer_205;
  reg        [31:0]   axi4Interface_fifoDataBuffer_206;
  reg        [31:0]   axi4Interface_fifoDataBuffer_207;
  reg        [31:0]   axi4Interface_fifoDataBuffer_208;
  reg        [31:0]   axi4Interface_fifoDataBuffer_209;
  reg        [31:0]   axi4Interface_fifoDataBuffer_210;
  reg        [31:0]   axi4Interface_fifoDataBuffer_211;
  reg        [31:0]   axi4Interface_fifoDataBuffer_212;
  reg        [31:0]   axi4Interface_fifoDataBuffer_213;
  reg        [31:0]   axi4Interface_fifoDataBuffer_214;
  reg        [31:0]   axi4Interface_fifoDataBuffer_215;
  reg        [31:0]   axi4Interface_fifoDataBuffer_216;
  reg        [31:0]   axi4Interface_fifoDataBuffer_217;
  reg        [31:0]   axi4Interface_fifoDataBuffer_218;
  reg        [31:0]   axi4Interface_fifoDataBuffer_219;
  reg        [31:0]   axi4Interface_fifoDataBuffer_220;
  reg        [31:0]   axi4Interface_fifoDataBuffer_221;
  reg        [31:0]   axi4Interface_fifoDataBuffer_222;
  reg        [31:0]   axi4Interface_fifoDataBuffer_223;
  reg        [31:0]   axi4Interface_fifoDataBuffer_224;
  reg        [31:0]   axi4Interface_fifoDataBuffer_225;
  reg        [31:0]   axi4Interface_fifoDataBuffer_226;
  reg        [31:0]   axi4Interface_fifoDataBuffer_227;
  reg        [31:0]   axi4Interface_fifoDataBuffer_228;
  reg        [31:0]   axi4Interface_fifoDataBuffer_229;
  reg        [31:0]   axi4Interface_fifoDataBuffer_230;
  reg        [31:0]   axi4Interface_fifoDataBuffer_231;
  reg        [31:0]   axi4Interface_fifoDataBuffer_232;
  reg        [31:0]   axi4Interface_fifoDataBuffer_233;
  reg        [31:0]   axi4Interface_fifoDataBuffer_234;
  reg        [31:0]   axi4Interface_fifoDataBuffer_235;
  reg        [31:0]   axi4Interface_fifoDataBuffer_236;
  reg        [31:0]   axi4Interface_fifoDataBuffer_237;
  reg        [31:0]   axi4Interface_fifoDataBuffer_238;
  reg        [31:0]   axi4Interface_fifoDataBuffer_239;
  reg        [31:0]   axi4Interface_fifoDataBuffer_240;
  reg        [31:0]   axi4Interface_fifoDataBuffer_241;
  reg        [31:0]   axi4Interface_fifoDataBuffer_242;
  reg        [31:0]   axi4Interface_fifoDataBuffer_243;
  reg        [31:0]   axi4Interface_fifoDataBuffer_244;
  reg        [31:0]   axi4Interface_fifoDataBuffer_245;
  reg        [31:0]   axi4Interface_fifoDataBuffer_246;
  reg        [31:0]   axi4Interface_fifoDataBuffer_247;
  reg        [31:0]   axi4Interface_fifoDataBuffer_248;
  reg        [31:0]   axi4Interface_fifoDataBuffer_249;
  reg        [31:0]   axi4Interface_fifoDataBuffer_250;
  reg        [31:0]   axi4Interface_fifoDataBuffer_251;
  reg        [31:0]   axi4Interface_fifoDataBuffer_252;
  reg        [31:0]   axi4Interface_fifoDataBuffer_253;
  reg        [31:0]   axi4Interface_fifoDataBuffer_254;
  reg        [31:0]   axi4Interface_fifoDataBuffer_255;
  wire                axi4Interface_stream_fire;
  wire       [255:0]  _zz_5;
  wire                when_Axi4WriteMaster_l55;
  reg        [31:0]   axi4Interface_address /* verilator public */ ;
  wire                axi4Interface_t_w_fire;
  wire       [1:0]    Axi4Incr_validSize;
  reg        [31:0]   Axi4Incr_result;
  wire       [19:0]   Axi4Incr_highCat;
  wire       [2:0]    Axi4Incr_sizeValue;
  wire       [11:0]   Axi4Incr_alignMask;
  wire       [11:0]   Axi4Incr_base;
  wire       [11:0]   Axi4Incr_baseIncr;
  reg        [1:0]    _zz_Axi4Incr_wrapCase;
  wire       [2:0]    Axi4Incr_wrapCase;
  reg                 axi4Interface_controlAwValid;
  reg                 axi4Interface_isTransferAfterReset;
  wire                axi4Interface_t_aw_fire;
  wire                when_Axi4WriteMaster_l92;
  reg        [31:0]   axi4Interface_initialAddress;
  wire                axi4Interface_t_w_fire_1;
  wire                when_Axi4WriteMaster_l141;
  reg                 axi4Interface_controlBReady;
  reg                 m_axi_wvalid_regNext;
  wire                when_Axi4WriteMaster_l156;
  wire                axi4Interface_t_b_fire;

  assign _zz__zz_m_axi_wdata_1_1 = _zz_m_axi_wdata;
  assign _zz__zz_m_axi_wdata_1 = {8'd0, _zz__zz_m_axi_wdata_1_1};
  assign _zz__zz_when_Axi4WriteMaster_l55_1_1 = _zz_when_Axi4WriteMaster_l55;
  assign _zz__zz_when_Axi4WriteMaster_l55_1 = {8'd0, _zz__zz_when_Axi4WriteMaster_l55_1_1};
  assign _zz__zz_5 = _zz_when_Axi4WriteMaster_l55_2[7:0];
  assign _zz_Axi4Incr_alignMask = {(2'b01 < Axi4Incr_validSize),(2'b00 < Axi4Incr_validSize)};
  assign _zz_Axi4Incr_base_1 = axi4Interface_address[11 : 0];
  assign _zz_Axi4Incr_base = _zz_Axi4Incr_base_1;
  assign _zz_Axi4Incr_baseIncr = {9'd0, Axi4Incr_sizeValue};
  assign _zz_Axi4Incr_wrapCase_1 = {1'd0, Axi4Incr_validSize};
  assign _zz_Axi4Incr_wrapCase_2 = {1'd0, _zz_Axi4Incr_wrapCase};
  assign _zz_m_axi_wdata_4 = _zz_m_axi_wdata_2[7:0];
  assign _zz_Axi4Incr_result_1 = Axi4Incr_base[11 : 1];
  assign _zz_Axi4Incr_result_2 = Axi4Incr_baseIncr[0 : 0];
  assign _zz_Axi4Incr_result_3 = Axi4Incr_base[11 : 2];
  assign _zz_Axi4Incr_result_4 = Axi4Incr_baseIncr[1 : 0];
  assign _zz_Axi4Incr_result_5 = Axi4Incr_base[11 : 3];
  assign _zz_Axi4Incr_result_6 = Axi4Incr_baseIncr[2 : 0];
  assign _zz_Axi4Incr_result_7 = Axi4Incr_base[11 : 4];
  assign _zz_Axi4Incr_result_8 = Axi4Incr_baseIncr[3 : 0];
  assign _zz_Axi4Incr_result_9 = Axi4Incr_base[11 : 5];
  assign _zz_Axi4Incr_result_10 = Axi4Incr_baseIncr[4 : 0];
  assign _zz_Axi4Incr_result_11 = Axi4Incr_base[11 : 6];
  assign _zz_Axi4Incr_result_12 = Axi4Incr_baseIncr[5 : 0];
  always @(*) begin
    case(Axi4Incr_wrapCase)
      3'b000 : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_1,_zz_Axi4Incr_result_2};
      end
      3'b001 : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_3,_zz_Axi4Incr_result_4};
      end
      3'b010 : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_5,_zz_Axi4Incr_result_6};
      end
      3'b011 : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_7,_zz_Axi4Incr_result_8};
      end
      3'b100 : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_9,_zz_Axi4Incr_result_10};
      end
      default : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_11,_zz_Axi4Incr_result_12};
      end
    endcase
  end

  always @(*) begin
    case(_zz_m_axi_wdata_4)
      8'b00000000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_0;
      end
      8'b00000001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_1;
      end
      8'b00000010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_2;
      end
      8'b00000011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_3;
      end
      8'b00000100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_4;
      end
      8'b00000101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_5;
      end
      8'b00000110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_6;
      end
      8'b00000111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_7;
      end
      8'b00001000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_8;
      end
      8'b00001001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_9;
      end
      8'b00001010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_10;
      end
      8'b00001011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_11;
      end
      8'b00001100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_12;
      end
      8'b00001101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_13;
      end
      8'b00001110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_14;
      end
      8'b00001111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_15;
      end
      8'b00010000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_16;
      end
      8'b00010001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_17;
      end
      8'b00010010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_18;
      end
      8'b00010011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_19;
      end
      8'b00010100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_20;
      end
      8'b00010101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_21;
      end
      8'b00010110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_22;
      end
      8'b00010111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_23;
      end
      8'b00011000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_24;
      end
      8'b00011001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_25;
      end
      8'b00011010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_26;
      end
      8'b00011011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_27;
      end
      8'b00011100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_28;
      end
      8'b00011101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_29;
      end
      8'b00011110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_30;
      end
      8'b00011111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_31;
      end
      8'b00100000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_32;
      end
      8'b00100001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_33;
      end
      8'b00100010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_34;
      end
      8'b00100011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_35;
      end
      8'b00100100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_36;
      end
      8'b00100101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_37;
      end
      8'b00100110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_38;
      end
      8'b00100111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_39;
      end
      8'b00101000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_40;
      end
      8'b00101001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_41;
      end
      8'b00101010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_42;
      end
      8'b00101011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_43;
      end
      8'b00101100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_44;
      end
      8'b00101101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_45;
      end
      8'b00101110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_46;
      end
      8'b00101111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_47;
      end
      8'b00110000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_48;
      end
      8'b00110001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_49;
      end
      8'b00110010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_50;
      end
      8'b00110011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_51;
      end
      8'b00110100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_52;
      end
      8'b00110101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_53;
      end
      8'b00110110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_54;
      end
      8'b00110111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_55;
      end
      8'b00111000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_56;
      end
      8'b00111001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_57;
      end
      8'b00111010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_58;
      end
      8'b00111011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_59;
      end
      8'b00111100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_60;
      end
      8'b00111101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_61;
      end
      8'b00111110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_62;
      end
      8'b00111111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_63;
      end
      8'b01000000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_64;
      end
      8'b01000001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_65;
      end
      8'b01000010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_66;
      end
      8'b01000011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_67;
      end
      8'b01000100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_68;
      end
      8'b01000101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_69;
      end
      8'b01000110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_70;
      end
      8'b01000111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_71;
      end
      8'b01001000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_72;
      end
      8'b01001001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_73;
      end
      8'b01001010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_74;
      end
      8'b01001011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_75;
      end
      8'b01001100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_76;
      end
      8'b01001101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_77;
      end
      8'b01001110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_78;
      end
      8'b01001111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_79;
      end
      8'b01010000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_80;
      end
      8'b01010001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_81;
      end
      8'b01010010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_82;
      end
      8'b01010011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_83;
      end
      8'b01010100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_84;
      end
      8'b01010101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_85;
      end
      8'b01010110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_86;
      end
      8'b01010111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_87;
      end
      8'b01011000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_88;
      end
      8'b01011001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_89;
      end
      8'b01011010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_90;
      end
      8'b01011011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_91;
      end
      8'b01011100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_92;
      end
      8'b01011101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_93;
      end
      8'b01011110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_94;
      end
      8'b01011111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_95;
      end
      8'b01100000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_96;
      end
      8'b01100001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_97;
      end
      8'b01100010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_98;
      end
      8'b01100011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_99;
      end
      8'b01100100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_100;
      end
      8'b01100101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_101;
      end
      8'b01100110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_102;
      end
      8'b01100111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_103;
      end
      8'b01101000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_104;
      end
      8'b01101001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_105;
      end
      8'b01101010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_106;
      end
      8'b01101011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_107;
      end
      8'b01101100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_108;
      end
      8'b01101101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_109;
      end
      8'b01101110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_110;
      end
      8'b01101111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_111;
      end
      8'b01110000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_112;
      end
      8'b01110001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_113;
      end
      8'b01110010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_114;
      end
      8'b01110011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_115;
      end
      8'b01110100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_116;
      end
      8'b01110101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_117;
      end
      8'b01110110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_118;
      end
      8'b01110111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_119;
      end
      8'b01111000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_120;
      end
      8'b01111001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_121;
      end
      8'b01111010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_122;
      end
      8'b01111011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_123;
      end
      8'b01111100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_124;
      end
      8'b01111101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_125;
      end
      8'b01111110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_126;
      end
      8'b01111111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_127;
      end
      8'b10000000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_128;
      end
      8'b10000001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_129;
      end
      8'b10000010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_130;
      end
      8'b10000011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_131;
      end
      8'b10000100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_132;
      end
      8'b10000101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_133;
      end
      8'b10000110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_134;
      end
      8'b10000111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_135;
      end
      8'b10001000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_136;
      end
      8'b10001001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_137;
      end
      8'b10001010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_138;
      end
      8'b10001011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_139;
      end
      8'b10001100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_140;
      end
      8'b10001101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_141;
      end
      8'b10001110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_142;
      end
      8'b10001111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_143;
      end
      8'b10010000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_144;
      end
      8'b10010001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_145;
      end
      8'b10010010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_146;
      end
      8'b10010011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_147;
      end
      8'b10010100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_148;
      end
      8'b10010101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_149;
      end
      8'b10010110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_150;
      end
      8'b10010111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_151;
      end
      8'b10011000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_152;
      end
      8'b10011001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_153;
      end
      8'b10011010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_154;
      end
      8'b10011011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_155;
      end
      8'b10011100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_156;
      end
      8'b10011101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_157;
      end
      8'b10011110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_158;
      end
      8'b10011111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_159;
      end
      8'b10100000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_160;
      end
      8'b10100001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_161;
      end
      8'b10100010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_162;
      end
      8'b10100011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_163;
      end
      8'b10100100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_164;
      end
      8'b10100101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_165;
      end
      8'b10100110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_166;
      end
      8'b10100111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_167;
      end
      8'b10101000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_168;
      end
      8'b10101001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_169;
      end
      8'b10101010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_170;
      end
      8'b10101011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_171;
      end
      8'b10101100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_172;
      end
      8'b10101101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_173;
      end
      8'b10101110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_174;
      end
      8'b10101111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_175;
      end
      8'b10110000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_176;
      end
      8'b10110001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_177;
      end
      8'b10110010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_178;
      end
      8'b10110011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_179;
      end
      8'b10110100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_180;
      end
      8'b10110101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_181;
      end
      8'b10110110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_182;
      end
      8'b10110111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_183;
      end
      8'b10111000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_184;
      end
      8'b10111001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_185;
      end
      8'b10111010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_186;
      end
      8'b10111011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_187;
      end
      8'b10111100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_188;
      end
      8'b10111101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_189;
      end
      8'b10111110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_190;
      end
      8'b10111111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_191;
      end
      8'b11000000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_192;
      end
      8'b11000001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_193;
      end
      8'b11000010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_194;
      end
      8'b11000011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_195;
      end
      8'b11000100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_196;
      end
      8'b11000101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_197;
      end
      8'b11000110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_198;
      end
      8'b11000111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_199;
      end
      8'b11001000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_200;
      end
      8'b11001001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_201;
      end
      8'b11001010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_202;
      end
      8'b11001011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_203;
      end
      8'b11001100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_204;
      end
      8'b11001101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_205;
      end
      8'b11001110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_206;
      end
      8'b11001111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_207;
      end
      8'b11010000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_208;
      end
      8'b11010001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_209;
      end
      8'b11010010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_210;
      end
      8'b11010011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_211;
      end
      8'b11010100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_212;
      end
      8'b11010101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_213;
      end
      8'b11010110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_214;
      end
      8'b11010111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_215;
      end
      8'b11011000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_216;
      end
      8'b11011001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_217;
      end
      8'b11011010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_218;
      end
      8'b11011011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_219;
      end
      8'b11011100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_220;
      end
      8'b11011101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_221;
      end
      8'b11011110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_222;
      end
      8'b11011111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_223;
      end
      8'b11100000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_224;
      end
      8'b11100001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_225;
      end
      8'b11100010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_226;
      end
      8'b11100011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_227;
      end
      8'b11100100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_228;
      end
      8'b11100101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_229;
      end
      8'b11100110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_230;
      end
      8'b11100111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_231;
      end
      8'b11101000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_232;
      end
      8'b11101001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_233;
      end
      8'b11101010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_234;
      end
      8'b11101011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_235;
      end
      8'b11101100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_236;
      end
      8'b11101101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_237;
      end
      8'b11101110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_238;
      end
      8'b11101111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_239;
      end
      8'b11110000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_240;
      end
      8'b11110001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_241;
      end
      8'b11110010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_242;
      end
      8'b11110011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_243;
      end
      8'b11110100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_244;
      end
      8'b11110101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_245;
      end
      8'b11110110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_246;
      end
      8'b11110111 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_247;
      end
      8'b11111000 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_248;
      end
      8'b11111001 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_249;
      end
      8'b11111010 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_250;
      end
      8'b11111011 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_251;
      end
      8'b11111100 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_252;
      end
      8'b11111101 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_253;
      end
      8'b11111110 : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_254;
      end
      default : begin
        _zz_m_axi_wdata_3 = axi4Interface_fifoDataBuffer_255;
      end
    endcase
  end

  always @(*) begin
    _zz_m_axi_wdata = 1'b0;
    if(axi4Interface_t_w_fire_1) begin
      _zz_m_axi_wdata = 1'b1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(_zz_when_Axi4WriteMaster_l92) begin
      _zz_1 = 1'b1;
    end
  end

  assign _zz_when_Axi4WriteMaster_l92 = (_zz_m_axi_wdata_2 == 9'h100);
  assign _zz_2 = (_zz_when_Axi4WriteMaster_l92 && _zz_m_axi_wdata);
  always @(*) begin
    if(_zz_2) begin
      _zz_m_axi_wdata_1 = 9'h0;
    end else begin
      _zz_m_axi_wdata_1 = (_zz_m_axi_wdata_2 + _zz__zz_m_axi_wdata_1);
    end
    if(_zz_1) begin
      _zz_m_axi_wdata_1 = 9'h0;
    end
  end

  always @(*) begin
    _zz_when_Axi4WriteMaster_l55 = 1'b0;
    if(axi4Interface_stream_fire) begin
      _zz_when_Axi4WriteMaster_l55 = 1'b1;
    end
  end

  always @(*) begin
    _zz_3 = 1'b0;
    if(_zz_when_Axi4WriteMaster_l92) begin
      _zz_3 = 1'b1;
    end
  end

  assign _zz_when_Axi4WriteMaster_l55_3 = (_zz_when_Axi4WriteMaster_l55_2 == 9'h100);
  assign _zz_4 = (_zz_when_Axi4WriteMaster_l55_3 && _zz_when_Axi4WriteMaster_l55);
  always @(*) begin
    if(_zz_4) begin
      _zz_when_Axi4WriteMaster_l55_1 = 9'h0;
    end else begin
      _zz_when_Axi4WriteMaster_l55_1 = (_zz_when_Axi4WriteMaster_l55_2 + _zz__zz_when_Axi4WriteMaster_l55_1);
    end
    if(_zz_3) begin
      _zz_when_Axi4WriteMaster_l55_1 = 9'h0;
    end
  end

  assign axi4Interface_stream_fire = (s_axis_valid && s_axis_ready);
  assign _zz_5 = ({255'd0,1'b1} <<< _zz__zz_5);
  always @(*) begin
    s_axis_ready = 1'b0;
    if(when_Axi4WriteMaster_l55) begin
      s_axis_ready = 1'b1;
    end
  end

  assign when_Axi4WriteMaster_l55 = (! _zz_when_Axi4WriteMaster_l55_3);
  assign axi4Interface_t_w_fire = (m_axi_wvalid && m_axi_wready);
  assign Axi4Incr_validSize = m_axi_awsize[1 : 0];
  assign Axi4Incr_highCat = axi4Interface_address[31 : 12];
  assign Axi4Incr_sizeValue = {(2'b10 == Axi4Incr_validSize),{(2'b01 == Axi4Incr_validSize),(2'b00 == Axi4Incr_validSize)}};
  assign Axi4Incr_alignMask = {10'd0, _zz_Axi4Incr_alignMask};
  assign Axi4Incr_base = (_zz_Axi4Incr_base & (~ Axi4Incr_alignMask));
  assign Axi4Incr_baseIncr = (Axi4Incr_base + _zz_Axi4Incr_baseIncr);
  always @(*) begin
    casez(m_axi_awlen)
      8'b????1??? : begin
        _zz_Axi4Incr_wrapCase = 2'b11;
      end
      8'b????01?? : begin
        _zz_Axi4Incr_wrapCase = 2'b10;
      end
      8'b????001? : begin
        _zz_Axi4Incr_wrapCase = 2'b01;
      end
      default : begin
        _zz_Axi4Incr_wrapCase = 2'b00;
      end
    endcase
  end

  assign Axi4Incr_wrapCase = (_zz_Axi4Incr_wrapCase_1 + _zz_Axi4Incr_wrapCase_2);
  always @(*) begin
    case(m_axi_awburst)
      2'b00 : begin
        Axi4Incr_result = axi4Interface_address;
      end
      2'b10 : begin
        Axi4Incr_result = {Axi4Incr_highCat,_zz_Axi4Incr_result};
      end
      default : begin
        Axi4Incr_result = {Axi4Incr_highCat,Axi4Incr_baseIncr};
      end
    endcase
  end

  assign axi4Interface_t_aw_fire = (m_axi_awvalid && m_axi_awready);
  assign when_Axi4WriteMaster_l92 = (_zz_when_Axi4WriteMaster_l92 || axi4Interface_isTransferAfterReset);
  assign m_axi_awvalid = axi4Interface_controlAwValid;
  always @(*) begin
    if(_zz_when_Axi4WriteMaster_l92) begin
      m_axi_awaddr = axi4Interface_address;
    end else begin
      m_axi_awaddr = axi4Interface_initialAddress;
    end
  end

  assign m_axi_awregion = 4'b0000;
  assign m_axi_awburst = 2'b01;
  assign m_axi_awlen = 8'hff;
  assign m_axi_awsize = 3'b010;
  assign m_axi_awcache = 4'b0000;
  assign m_axi_awqos = 4'b0000;
  assign m_axi_awprot = 3'b000;
  always @(*) begin
    m_axi_wdata = 32'h0;
    if(m_axi_wvalid) begin
      m_axi_wdata = _zz_m_axi_wdata_3;
    end
  end

  assign axi4Interface_t_w_fire_1 = (m_axi_wvalid && m_axi_wready);
  always @(*) begin
    m_axi_wvalid = 1'b0;
    if(when_Axi4WriteMaster_l141) begin
      m_axi_wvalid = 1'b1;
    end
  end

  assign when_Axi4WriteMaster_l141 = (((9'h0 < _zz_when_Axi4WriteMaster_l55_2) && (_zz_m_axi_wdata_2 < _zz_when_Axi4WriteMaster_l55_2)) && (! _zz_when_Axi4WriteMaster_l92));
  assign m_axi_wstrb = 4'b1111;
  assign m_axi_wlast = (_zz_m_axi_wdata_2 == 9'h0ff);
  assign when_Axi4WriteMaster_l156 = (m_axi_wvalid && (! m_axi_wvalid_regNext));
  assign axi4Interface_t_b_fire = (m_axi_bvalid && m_axi_bready);
  assign m_axi_bready = axi4Interface_controlBReady;
  assign m_axi_araddr = 32'h0;
  assign m_axi_arregion = 4'b0000;
  assign m_axi_arburst = 2'b01;
  assign m_axi_arlen = 8'hff;
  assign m_axi_arsize = 3'b100;
  assign m_axi_arcache = 4'b0000;
  assign m_axi_arqos = 4'b0000;
  assign m_axi_arprot = 3'b000;
  assign m_axi_arvalid = 1'b0;
  assign m_axi_rready = 1'b0;
  always @(posedge aclk or posedge aresetn) begin
    if(aresetn) begin
      _zz_m_axi_wdata_2 <= 9'h0;
      _zz_when_Axi4WriteMaster_l55_2 <= 9'h0;
      axi4Interface_fifoDataBuffer_0 <= 32'h0;
      axi4Interface_fifoDataBuffer_1 <= 32'h0;
      axi4Interface_fifoDataBuffer_2 <= 32'h0;
      axi4Interface_fifoDataBuffer_3 <= 32'h0;
      axi4Interface_fifoDataBuffer_4 <= 32'h0;
      axi4Interface_fifoDataBuffer_5 <= 32'h0;
      axi4Interface_fifoDataBuffer_6 <= 32'h0;
      axi4Interface_fifoDataBuffer_7 <= 32'h0;
      axi4Interface_fifoDataBuffer_8 <= 32'h0;
      axi4Interface_fifoDataBuffer_9 <= 32'h0;
      axi4Interface_fifoDataBuffer_10 <= 32'h0;
      axi4Interface_fifoDataBuffer_11 <= 32'h0;
      axi4Interface_fifoDataBuffer_12 <= 32'h0;
      axi4Interface_fifoDataBuffer_13 <= 32'h0;
      axi4Interface_fifoDataBuffer_14 <= 32'h0;
      axi4Interface_fifoDataBuffer_15 <= 32'h0;
      axi4Interface_fifoDataBuffer_16 <= 32'h0;
      axi4Interface_fifoDataBuffer_17 <= 32'h0;
      axi4Interface_fifoDataBuffer_18 <= 32'h0;
      axi4Interface_fifoDataBuffer_19 <= 32'h0;
      axi4Interface_fifoDataBuffer_20 <= 32'h0;
      axi4Interface_fifoDataBuffer_21 <= 32'h0;
      axi4Interface_fifoDataBuffer_22 <= 32'h0;
      axi4Interface_fifoDataBuffer_23 <= 32'h0;
      axi4Interface_fifoDataBuffer_24 <= 32'h0;
      axi4Interface_fifoDataBuffer_25 <= 32'h0;
      axi4Interface_fifoDataBuffer_26 <= 32'h0;
      axi4Interface_fifoDataBuffer_27 <= 32'h0;
      axi4Interface_fifoDataBuffer_28 <= 32'h0;
      axi4Interface_fifoDataBuffer_29 <= 32'h0;
      axi4Interface_fifoDataBuffer_30 <= 32'h0;
      axi4Interface_fifoDataBuffer_31 <= 32'h0;
      axi4Interface_fifoDataBuffer_32 <= 32'h0;
      axi4Interface_fifoDataBuffer_33 <= 32'h0;
      axi4Interface_fifoDataBuffer_34 <= 32'h0;
      axi4Interface_fifoDataBuffer_35 <= 32'h0;
      axi4Interface_fifoDataBuffer_36 <= 32'h0;
      axi4Interface_fifoDataBuffer_37 <= 32'h0;
      axi4Interface_fifoDataBuffer_38 <= 32'h0;
      axi4Interface_fifoDataBuffer_39 <= 32'h0;
      axi4Interface_fifoDataBuffer_40 <= 32'h0;
      axi4Interface_fifoDataBuffer_41 <= 32'h0;
      axi4Interface_fifoDataBuffer_42 <= 32'h0;
      axi4Interface_fifoDataBuffer_43 <= 32'h0;
      axi4Interface_fifoDataBuffer_44 <= 32'h0;
      axi4Interface_fifoDataBuffer_45 <= 32'h0;
      axi4Interface_fifoDataBuffer_46 <= 32'h0;
      axi4Interface_fifoDataBuffer_47 <= 32'h0;
      axi4Interface_fifoDataBuffer_48 <= 32'h0;
      axi4Interface_fifoDataBuffer_49 <= 32'h0;
      axi4Interface_fifoDataBuffer_50 <= 32'h0;
      axi4Interface_fifoDataBuffer_51 <= 32'h0;
      axi4Interface_fifoDataBuffer_52 <= 32'h0;
      axi4Interface_fifoDataBuffer_53 <= 32'h0;
      axi4Interface_fifoDataBuffer_54 <= 32'h0;
      axi4Interface_fifoDataBuffer_55 <= 32'h0;
      axi4Interface_fifoDataBuffer_56 <= 32'h0;
      axi4Interface_fifoDataBuffer_57 <= 32'h0;
      axi4Interface_fifoDataBuffer_58 <= 32'h0;
      axi4Interface_fifoDataBuffer_59 <= 32'h0;
      axi4Interface_fifoDataBuffer_60 <= 32'h0;
      axi4Interface_fifoDataBuffer_61 <= 32'h0;
      axi4Interface_fifoDataBuffer_62 <= 32'h0;
      axi4Interface_fifoDataBuffer_63 <= 32'h0;
      axi4Interface_fifoDataBuffer_64 <= 32'h0;
      axi4Interface_fifoDataBuffer_65 <= 32'h0;
      axi4Interface_fifoDataBuffer_66 <= 32'h0;
      axi4Interface_fifoDataBuffer_67 <= 32'h0;
      axi4Interface_fifoDataBuffer_68 <= 32'h0;
      axi4Interface_fifoDataBuffer_69 <= 32'h0;
      axi4Interface_fifoDataBuffer_70 <= 32'h0;
      axi4Interface_fifoDataBuffer_71 <= 32'h0;
      axi4Interface_fifoDataBuffer_72 <= 32'h0;
      axi4Interface_fifoDataBuffer_73 <= 32'h0;
      axi4Interface_fifoDataBuffer_74 <= 32'h0;
      axi4Interface_fifoDataBuffer_75 <= 32'h0;
      axi4Interface_fifoDataBuffer_76 <= 32'h0;
      axi4Interface_fifoDataBuffer_77 <= 32'h0;
      axi4Interface_fifoDataBuffer_78 <= 32'h0;
      axi4Interface_fifoDataBuffer_79 <= 32'h0;
      axi4Interface_fifoDataBuffer_80 <= 32'h0;
      axi4Interface_fifoDataBuffer_81 <= 32'h0;
      axi4Interface_fifoDataBuffer_82 <= 32'h0;
      axi4Interface_fifoDataBuffer_83 <= 32'h0;
      axi4Interface_fifoDataBuffer_84 <= 32'h0;
      axi4Interface_fifoDataBuffer_85 <= 32'h0;
      axi4Interface_fifoDataBuffer_86 <= 32'h0;
      axi4Interface_fifoDataBuffer_87 <= 32'h0;
      axi4Interface_fifoDataBuffer_88 <= 32'h0;
      axi4Interface_fifoDataBuffer_89 <= 32'h0;
      axi4Interface_fifoDataBuffer_90 <= 32'h0;
      axi4Interface_fifoDataBuffer_91 <= 32'h0;
      axi4Interface_fifoDataBuffer_92 <= 32'h0;
      axi4Interface_fifoDataBuffer_93 <= 32'h0;
      axi4Interface_fifoDataBuffer_94 <= 32'h0;
      axi4Interface_fifoDataBuffer_95 <= 32'h0;
      axi4Interface_fifoDataBuffer_96 <= 32'h0;
      axi4Interface_fifoDataBuffer_97 <= 32'h0;
      axi4Interface_fifoDataBuffer_98 <= 32'h0;
      axi4Interface_fifoDataBuffer_99 <= 32'h0;
      axi4Interface_fifoDataBuffer_100 <= 32'h0;
      axi4Interface_fifoDataBuffer_101 <= 32'h0;
      axi4Interface_fifoDataBuffer_102 <= 32'h0;
      axi4Interface_fifoDataBuffer_103 <= 32'h0;
      axi4Interface_fifoDataBuffer_104 <= 32'h0;
      axi4Interface_fifoDataBuffer_105 <= 32'h0;
      axi4Interface_fifoDataBuffer_106 <= 32'h0;
      axi4Interface_fifoDataBuffer_107 <= 32'h0;
      axi4Interface_fifoDataBuffer_108 <= 32'h0;
      axi4Interface_fifoDataBuffer_109 <= 32'h0;
      axi4Interface_fifoDataBuffer_110 <= 32'h0;
      axi4Interface_fifoDataBuffer_111 <= 32'h0;
      axi4Interface_fifoDataBuffer_112 <= 32'h0;
      axi4Interface_fifoDataBuffer_113 <= 32'h0;
      axi4Interface_fifoDataBuffer_114 <= 32'h0;
      axi4Interface_fifoDataBuffer_115 <= 32'h0;
      axi4Interface_fifoDataBuffer_116 <= 32'h0;
      axi4Interface_fifoDataBuffer_117 <= 32'h0;
      axi4Interface_fifoDataBuffer_118 <= 32'h0;
      axi4Interface_fifoDataBuffer_119 <= 32'h0;
      axi4Interface_fifoDataBuffer_120 <= 32'h0;
      axi4Interface_fifoDataBuffer_121 <= 32'h0;
      axi4Interface_fifoDataBuffer_122 <= 32'h0;
      axi4Interface_fifoDataBuffer_123 <= 32'h0;
      axi4Interface_fifoDataBuffer_124 <= 32'h0;
      axi4Interface_fifoDataBuffer_125 <= 32'h0;
      axi4Interface_fifoDataBuffer_126 <= 32'h0;
      axi4Interface_fifoDataBuffer_127 <= 32'h0;
      axi4Interface_fifoDataBuffer_128 <= 32'h0;
      axi4Interface_fifoDataBuffer_129 <= 32'h0;
      axi4Interface_fifoDataBuffer_130 <= 32'h0;
      axi4Interface_fifoDataBuffer_131 <= 32'h0;
      axi4Interface_fifoDataBuffer_132 <= 32'h0;
      axi4Interface_fifoDataBuffer_133 <= 32'h0;
      axi4Interface_fifoDataBuffer_134 <= 32'h0;
      axi4Interface_fifoDataBuffer_135 <= 32'h0;
      axi4Interface_fifoDataBuffer_136 <= 32'h0;
      axi4Interface_fifoDataBuffer_137 <= 32'h0;
      axi4Interface_fifoDataBuffer_138 <= 32'h0;
      axi4Interface_fifoDataBuffer_139 <= 32'h0;
      axi4Interface_fifoDataBuffer_140 <= 32'h0;
      axi4Interface_fifoDataBuffer_141 <= 32'h0;
      axi4Interface_fifoDataBuffer_142 <= 32'h0;
      axi4Interface_fifoDataBuffer_143 <= 32'h0;
      axi4Interface_fifoDataBuffer_144 <= 32'h0;
      axi4Interface_fifoDataBuffer_145 <= 32'h0;
      axi4Interface_fifoDataBuffer_146 <= 32'h0;
      axi4Interface_fifoDataBuffer_147 <= 32'h0;
      axi4Interface_fifoDataBuffer_148 <= 32'h0;
      axi4Interface_fifoDataBuffer_149 <= 32'h0;
      axi4Interface_fifoDataBuffer_150 <= 32'h0;
      axi4Interface_fifoDataBuffer_151 <= 32'h0;
      axi4Interface_fifoDataBuffer_152 <= 32'h0;
      axi4Interface_fifoDataBuffer_153 <= 32'h0;
      axi4Interface_fifoDataBuffer_154 <= 32'h0;
      axi4Interface_fifoDataBuffer_155 <= 32'h0;
      axi4Interface_fifoDataBuffer_156 <= 32'h0;
      axi4Interface_fifoDataBuffer_157 <= 32'h0;
      axi4Interface_fifoDataBuffer_158 <= 32'h0;
      axi4Interface_fifoDataBuffer_159 <= 32'h0;
      axi4Interface_fifoDataBuffer_160 <= 32'h0;
      axi4Interface_fifoDataBuffer_161 <= 32'h0;
      axi4Interface_fifoDataBuffer_162 <= 32'h0;
      axi4Interface_fifoDataBuffer_163 <= 32'h0;
      axi4Interface_fifoDataBuffer_164 <= 32'h0;
      axi4Interface_fifoDataBuffer_165 <= 32'h0;
      axi4Interface_fifoDataBuffer_166 <= 32'h0;
      axi4Interface_fifoDataBuffer_167 <= 32'h0;
      axi4Interface_fifoDataBuffer_168 <= 32'h0;
      axi4Interface_fifoDataBuffer_169 <= 32'h0;
      axi4Interface_fifoDataBuffer_170 <= 32'h0;
      axi4Interface_fifoDataBuffer_171 <= 32'h0;
      axi4Interface_fifoDataBuffer_172 <= 32'h0;
      axi4Interface_fifoDataBuffer_173 <= 32'h0;
      axi4Interface_fifoDataBuffer_174 <= 32'h0;
      axi4Interface_fifoDataBuffer_175 <= 32'h0;
      axi4Interface_fifoDataBuffer_176 <= 32'h0;
      axi4Interface_fifoDataBuffer_177 <= 32'h0;
      axi4Interface_fifoDataBuffer_178 <= 32'h0;
      axi4Interface_fifoDataBuffer_179 <= 32'h0;
      axi4Interface_fifoDataBuffer_180 <= 32'h0;
      axi4Interface_fifoDataBuffer_181 <= 32'h0;
      axi4Interface_fifoDataBuffer_182 <= 32'h0;
      axi4Interface_fifoDataBuffer_183 <= 32'h0;
      axi4Interface_fifoDataBuffer_184 <= 32'h0;
      axi4Interface_fifoDataBuffer_185 <= 32'h0;
      axi4Interface_fifoDataBuffer_186 <= 32'h0;
      axi4Interface_fifoDataBuffer_187 <= 32'h0;
      axi4Interface_fifoDataBuffer_188 <= 32'h0;
      axi4Interface_fifoDataBuffer_189 <= 32'h0;
      axi4Interface_fifoDataBuffer_190 <= 32'h0;
      axi4Interface_fifoDataBuffer_191 <= 32'h0;
      axi4Interface_fifoDataBuffer_192 <= 32'h0;
      axi4Interface_fifoDataBuffer_193 <= 32'h0;
      axi4Interface_fifoDataBuffer_194 <= 32'h0;
      axi4Interface_fifoDataBuffer_195 <= 32'h0;
      axi4Interface_fifoDataBuffer_196 <= 32'h0;
      axi4Interface_fifoDataBuffer_197 <= 32'h0;
      axi4Interface_fifoDataBuffer_198 <= 32'h0;
      axi4Interface_fifoDataBuffer_199 <= 32'h0;
      axi4Interface_fifoDataBuffer_200 <= 32'h0;
      axi4Interface_fifoDataBuffer_201 <= 32'h0;
      axi4Interface_fifoDataBuffer_202 <= 32'h0;
      axi4Interface_fifoDataBuffer_203 <= 32'h0;
      axi4Interface_fifoDataBuffer_204 <= 32'h0;
      axi4Interface_fifoDataBuffer_205 <= 32'h0;
      axi4Interface_fifoDataBuffer_206 <= 32'h0;
      axi4Interface_fifoDataBuffer_207 <= 32'h0;
      axi4Interface_fifoDataBuffer_208 <= 32'h0;
      axi4Interface_fifoDataBuffer_209 <= 32'h0;
      axi4Interface_fifoDataBuffer_210 <= 32'h0;
      axi4Interface_fifoDataBuffer_211 <= 32'h0;
      axi4Interface_fifoDataBuffer_212 <= 32'h0;
      axi4Interface_fifoDataBuffer_213 <= 32'h0;
      axi4Interface_fifoDataBuffer_214 <= 32'h0;
      axi4Interface_fifoDataBuffer_215 <= 32'h0;
      axi4Interface_fifoDataBuffer_216 <= 32'h0;
      axi4Interface_fifoDataBuffer_217 <= 32'h0;
      axi4Interface_fifoDataBuffer_218 <= 32'h0;
      axi4Interface_fifoDataBuffer_219 <= 32'h0;
      axi4Interface_fifoDataBuffer_220 <= 32'h0;
      axi4Interface_fifoDataBuffer_221 <= 32'h0;
      axi4Interface_fifoDataBuffer_222 <= 32'h0;
      axi4Interface_fifoDataBuffer_223 <= 32'h0;
      axi4Interface_fifoDataBuffer_224 <= 32'h0;
      axi4Interface_fifoDataBuffer_225 <= 32'h0;
      axi4Interface_fifoDataBuffer_226 <= 32'h0;
      axi4Interface_fifoDataBuffer_227 <= 32'h0;
      axi4Interface_fifoDataBuffer_228 <= 32'h0;
      axi4Interface_fifoDataBuffer_229 <= 32'h0;
      axi4Interface_fifoDataBuffer_230 <= 32'h0;
      axi4Interface_fifoDataBuffer_231 <= 32'h0;
      axi4Interface_fifoDataBuffer_232 <= 32'h0;
      axi4Interface_fifoDataBuffer_233 <= 32'h0;
      axi4Interface_fifoDataBuffer_234 <= 32'h0;
      axi4Interface_fifoDataBuffer_235 <= 32'h0;
      axi4Interface_fifoDataBuffer_236 <= 32'h0;
      axi4Interface_fifoDataBuffer_237 <= 32'h0;
      axi4Interface_fifoDataBuffer_238 <= 32'h0;
      axi4Interface_fifoDataBuffer_239 <= 32'h0;
      axi4Interface_fifoDataBuffer_240 <= 32'h0;
      axi4Interface_fifoDataBuffer_241 <= 32'h0;
      axi4Interface_fifoDataBuffer_242 <= 32'h0;
      axi4Interface_fifoDataBuffer_243 <= 32'h0;
      axi4Interface_fifoDataBuffer_244 <= 32'h0;
      axi4Interface_fifoDataBuffer_245 <= 32'h0;
      axi4Interface_fifoDataBuffer_246 <= 32'h0;
      axi4Interface_fifoDataBuffer_247 <= 32'h0;
      axi4Interface_fifoDataBuffer_248 <= 32'h0;
      axi4Interface_fifoDataBuffer_249 <= 32'h0;
      axi4Interface_fifoDataBuffer_250 <= 32'h0;
      axi4Interface_fifoDataBuffer_251 <= 32'h0;
      axi4Interface_fifoDataBuffer_252 <= 32'h0;
      axi4Interface_fifoDataBuffer_253 <= 32'h0;
      axi4Interface_fifoDataBuffer_254 <= 32'h0;
      axi4Interface_fifoDataBuffer_255 <= 32'h0;
      axi4Interface_address <= 32'h0;
      axi4Interface_controlAwValid <= 1'b0;
      axi4Interface_isTransferAfterReset <= 1'b1;
      axi4Interface_initialAddress <= 32'h0;
      axi4Interface_controlBReady <= 1'b0;
    end else begin
      _zz_m_axi_wdata_2 <= _zz_m_axi_wdata_1;
      _zz_when_Axi4WriteMaster_l55_2 <= _zz_when_Axi4WriteMaster_l55_1;
      if(axi4Interface_stream_fire) begin
        if(_zz_5[0]) begin
          axi4Interface_fifoDataBuffer_0 <= s_axis_payload;
        end
        if(_zz_5[1]) begin
          axi4Interface_fifoDataBuffer_1 <= s_axis_payload;
        end
        if(_zz_5[2]) begin
          axi4Interface_fifoDataBuffer_2 <= s_axis_payload;
        end
        if(_zz_5[3]) begin
          axi4Interface_fifoDataBuffer_3 <= s_axis_payload;
        end
        if(_zz_5[4]) begin
          axi4Interface_fifoDataBuffer_4 <= s_axis_payload;
        end
        if(_zz_5[5]) begin
          axi4Interface_fifoDataBuffer_5 <= s_axis_payload;
        end
        if(_zz_5[6]) begin
          axi4Interface_fifoDataBuffer_6 <= s_axis_payload;
        end
        if(_zz_5[7]) begin
          axi4Interface_fifoDataBuffer_7 <= s_axis_payload;
        end
        if(_zz_5[8]) begin
          axi4Interface_fifoDataBuffer_8 <= s_axis_payload;
        end
        if(_zz_5[9]) begin
          axi4Interface_fifoDataBuffer_9 <= s_axis_payload;
        end
        if(_zz_5[10]) begin
          axi4Interface_fifoDataBuffer_10 <= s_axis_payload;
        end
        if(_zz_5[11]) begin
          axi4Interface_fifoDataBuffer_11 <= s_axis_payload;
        end
        if(_zz_5[12]) begin
          axi4Interface_fifoDataBuffer_12 <= s_axis_payload;
        end
        if(_zz_5[13]) begin
          axi4Interface_fifoDataBuffer_13 <= s_axis_payload;
        end
        if(_zz_5[14]) begin
          axi4Interface_fifoDataBuffer_14 <= s_axis_payload;
        end
        if(_zz_5[15]) begin
          axi4Interface_fifoDataBuffer_15 <= s_axis_payload;
        end
        if(_zz_5[16]) begin
          axi4Interface_fifoDataBuffer_16 <= s_axis_payload;
        end
        if(_zz_5[17]) begin
          axi4Interface_fifoDataBuffer_17 <= s_axis_payload;
        end
        if(_zz_5[18]) begin
          axi4Interface_fifoDataBuffer_18 <= s_axis_payload;
        end
        if(_zz_5[19]) begin
          axi4Interface_fifoDataBuffer_19 <= s_axis_payload;
        end
        if(_zz_5[20]) begin
          axi4Interface_fifoDataBuffer_20 <= s_axis_payload;
        end
        if(_zz_5[21]) begin
          axi4Interface_fifoDataBuffer_21 <= s_axis_payload;
        end
        if(_zz_5[22]) begin
          axi4Interface_fifoDataBuffer_22 <= s_axis_payload;
        end
        if(_zz_5[23]) begin
          axi4Interface_fifoDataBuffer_23 <= s_axis_payload;
        end
        if(_zz_5[24]) begin
          axi4Interface_fifoDataBuffer_24 <= s_axis_payload;
        end
        if(_zz_5[25]) begin
          axi4Interface_fifoDataBuffer_25 <= s_axis_payload;
        end
        if(_zz_5[26]) begin
          axi4Interface_fifoDataBuffer_26 <= s_axis_payload;
        end
        if(_zz_5[27]) begin
          axi4Interface_fifoDataBuffer_27 <= s_axis_payload;
        end
        if(_zz_5[28]) begin
          axi4Interface_fifoDataBuffer_28 <= s_axis_payload;
        end
        if(_zz_5[29]) begin
          axi4Interface_fifoDataBuffer_29 <= s_axis_payload;
        end
        if(_zz_5[30]) begin
          axi4Interface_fifoDataBuffer_30 <= s_axis_payload;
        end
        if(_zz_5[31]) begin
          axi4Interface_fifoDataBuffer_31 <= s_axis_payload;
        end
        if(_zz_5[32]) begin
          axi4Interface_fifoDataBuffer_32 <= s_axis_payload;
        end
        if(_zz_5[33]) begin
          axi4Interface_fifoDataBuffer_33 <= s_axis_payload;
        end
        if(_zz_5[34]) begin
          axi4Interface_fifoDataBuffer_34 <= s_axis_payload;
        end
        if(_zz_5[35]) begin
          axi4Interface_fifoDataBuffer_35 <= s_axis_payload;
        end
        if(_zz_5[36]) begin
          axi4Interface_fifoDataBuffer_36 <= s_axis_payload;
        end
        if(_zz_5[37]) begin
          axi4Interface_fifoDataBuffer_37 <= s_axis_payload;
        end
        if(_zz_5[38]) begin
          axi4Interface_fifoDataBuffer_38 <= s_axis_payload;
        end
        if(_zz_5[39]) begin
          axi4Interface_fifoDataBuffer_39 <= s_axis_payload;
        end
        if(_zz_5[40]) begin
          axi4Interface_fifoDataBuffer_40 <= s_axis_payload;
        end
        if(_zz_5[41]) begin
          axi4Interface_fifoDataBuffer_41 <= s_axis_payload;
        end
        if(_zz_5[42]) begin
          axi4Interface_fifoDataBuffer_42 <= s_axis_payload;
        end
        if(_zz_5[43]) begin
          axi4Interface_fifoDataBuffer_43 <= s_axis_payload;
        end
        if(_zz_5[44]) begin
          axi4Interface_fifoDataBuffer_44 <= s_axis_payload;
        end
        if(_zz_5[45]) begin
          axi4Interface_fifoDataBuffer_45 <= s_axis_payload;
        end
        if(_zz_5[46]) begin
          axi4Interface_fifoDataBuffer_46 <= s_axis_payload;
        end
        if(_zz_5[47]) begin
          axi4Interface_fifoDataBuffer_47 <= s_axis_payload;
        end
        if(_zz_5[48]) begin
          axi4Interface_fifoDataBuffer_48 <= s_axis_payload;
        end
        if(_zz_5[49]) begin
          axi4Interface_fifoDataBuffer_49 <= s_axis_payload;
        end
        if(_zz_5[50]) begin
          axi4Interface_fifoDataBuffer_50 <= s_axis_payload;
        end
        if(_zz_5[51]) begin
          axi4Interface_fifoDataBuffer_51 <= s_axis_payload;
        end
        if(_zz_5[52]) begin
          axi4Interface_fifoDataBuffer_52 <= s_axis_payload;
        end
        if(_zz_5[53]) begin
          axi4Interface_fifoDataBuffer_53 <= s_axis_payload;
        end
        if(_zz_5[54]) begin
          axi4Interface_fifoDataBuffer_54 <= s_axis_payload;
        end
        if(_zz_5[55]) begin
          axi4Interface_fifoDataBuffer_55 <= s_axis_payload;
        end
        if(_zz_5[56]) begin
          axi4Interface_fifoDataBuffer_56 <= s_axis_payload;
        end
        if(_zz_5[57]) begin
          axi4Interface_fifoDataBuffer_57 <= s_axis_payload;
        end
        if(_zz_5[58]) begin
          axi4Interface_fifoDataBuffer_58 <= s_axis_payload;
        end
        if(_zz_5[59]) begin
          axi4Interface_fifoDataBuffer_59 <= s_axis_payload;
        end
        if(_zz_5[60]) begin
          axi4Interface_fifoDataBuffer_60 <= s_axis_payload;
        end
        if(_zz_5[61]) begin
          axi4Interface_fifoDataBuffer_61 <= s_axis_payload;
        end
        if(_zz_5[62]) begin
          axi4Interface_fifoDataBuffer_62 <= s_axis_payload;
        end
        if(_zz_5[63]) begin
          axi4Interface_fifoDataBuffer_63 <= s_axis_payload;
        end
        if(_zz_5[64]) begin
          axi4Interface_fifoDataBuffer_64 <= s_axis_payload;
        end
        if(_zz_5[65]) begin
          axi4Interface_fifoDataBuffer_65 <= s_axis_payload;
        end
        if(_zz_5[66]) begin
          axi4Interface_fifoDataBuffer_66 <= s_axis_payload;
        end
        if(_zz_5[67]) begin
          axi4Interface_fifoDataBuffer_67 <= s_axis_payload;
        end
        if(_zz_5[68]) begin
          axi4Interface_fifoDataBuffer_68 <= s_axis_payload;
        end
        if(_zz_5[69]) begin
          axi4Interface_fifoDataBuffer_69 <= s_axis_payload;
        end
        if(_zz_5[70]) begin
          axi4Interface_fifoDataBuffer_70 <= s_axis_payload;
        end
        if(_zz_5[71]) begin
          axi4Interface_fifoDataBuffer_71 <= s_axis_payload;
        end
        if(_zz_5[72]) begin
          axi4Interface_fifoDataBuffer_72 <= s_axis_payload;
        end
        if(_zz_5[73]) begin
          axi4Interface_fifoDataBuffer_73 <= s_axis_payload;
        end
        if(_zz_5[74]) begin
          axi4Interface_fifoDataBuffer_74 <= s_axis_payload;
        end
        if(_zz_5[75]) begin
          axi4Interface_fifoDataBuffer_75 <= s_axis_payload;
        end
        if(_zz_5[76]) begin
          axi4Interface_fifoDataBuffer_76 <= s_axis_payload;
        end
        if(_zz_5[77]) begin
          axi4Interface_fifoDataBuffer_77 <= s_axis_payload;
        end
        if(_zz_5[78]) begin
          axi4Interface_fifoDataBuffer_78 <= s_axis_payload;
        end
        if(_zz_5[79]) begin
          axi4Interface_fifoDataBuffer_79 <= s_axis_payload;
        end
        if(_zz_5[80]) begin
          axi4Interface_fifoDataBuffer_80 <= s_axis_payload;
        end
        if(_zz_5[81]) begin
          axi4Interface_fifoDataBuffer_81 <= s_axis_payload;
        end
        if(_zz_5[82]) begin
          axi4Interface_fifoDataBuffer_82 <= s_axis_payload;
        end
        if(_zz_5[83]) begin
          axi4Interface_fifoDataBuffer_83 <= s_axis_payload;
        end
        if(_zz_5[84]) begin
          axi4Interface_fifoDataBuffer_84 <= s_axis_payload;
        end
        if(_zz_5[85]) begin
          axi4Interface_fifoDataBuffer_85 <= s_axis_payload;
        end
        if(_zz_5[86]) begin
          axi4Interface_fifoDataBuffer_86 <= s_axis_payload;
        end
        if(_zz_5[87]) begin
          axi4Interface_fifoDataBuffer_87 <= s_axis_payload;
        end
        if(_zz_5[88]) begin
          axi4Interface_fifoDataBuffer_88 <= s_axis_payload;
        end
        if(_zz_5[89]) begin
          axi4Interface_fifoDataBuffer_89 <= s_axis_payload;
        end
        if(_zz_5[90]) begin
          axi4Interface_fifoDataBuffer_90 <= s_axis_payload;
        end
        if(_zz_5[91]) begin
          axi4Interface_fifoDataBuffer_91 <= s_axis_payload;
        end
        if(_zz_5[92]) begin
          axi4Interface_fifoDataBuffer_92 <= s_axis_payload;
        end
        if(_zz_5[93]) begin
          axi4Interface_fifoDataBuffer_93 <= s_axis_payload;
        end
        if(_zz_5[94]) begin
          axi4Interface_fifoDataBuffer_94 <= s_axis_payload;
        end
        if(_zz_5[95]) begin
          axi4Interface_fifoDataBuffer_95 <= s_axis_payload;
        end
        if(_zz_5[96]) begin
          axi4Interface_fifoDataBuffer_96 <= s_axis_payload;
        end
        if(_zz_5[97]) begin
          axi4Interface_fifoDataBuffer_97 <= s_axis_payload;
        end
        if(_zz_5[98]) begin
          axi4Interface_fifoDataBuffer_98 <= s_axis_payload;
        end
        if(_zz_5[99]) begin
          axi4Interface_fifoDataBuffer_99 <= s_axis_payload;
        end
        if(_zz_5[100]) begin
          axi4Interface_fifoDataBuffer_100 <= s_axis_payload;
        end
        if(_zz_5[101]) begin
          axi4Interface_fifoDataBuffer_101 <= s_axis_payload;
        end
        if(_zz_5[102]) begin
          axi4Interface_fifoDataBuffer_102 <= s_axis_payload;
        end
        if(_zz_5[103]) begin
          axi4Interface_fifoDataBuffer_103 <= s_axis_payload;
        end
        if(_zz_5[104]) begin
          axi4Interface_fifoDataBuffer_104 <= s_axis_payload;
        end
        if(_zz_5[105]) begin
          axi4Interface_fifoDataBuffer_105 <= s_axis_payload;
        end
        if(_zz_5[106]) begin
          axi4Interface_fifoDataBuffer_106 <= s_axis_payload;
        end
        if(_zz_5[107]) begin
          axi4Interface_fifoDataBuffer_107 <= s_axis_payload;
        end
        if(_zz_5[108]) begin
          axi4Interface_fifoDataBuffer_108 <= s_axis_payload;
        end
        if(_zz_5[109]) begin
          axi4Interface_fifoDataBuffer_109 <= s_axis_payload;
        end
        if(_zz_5[110]) begin
          axi4Interface_fifoDataBuffer_110 <= s_axis_payload;
        end
        if(_zz_5[111]) begin
          axi4Interface_fifoDataBuffer_111 <= s_axis_payload;
        end
        if(_zz_5[112]) begin
          axi4Interface_fifoDataBuffer_112 <= s_axis_payload;
        end
        if(_zz_5[113]) begin
          axi4Interface_fifoDataBuffer_113 <= s_axis_payload;
        end
        if(_zz_5[114]) begin
          axi4Interface_fifoDataBuffer_114 <= s_axis_payload;
        end
        if(_zz_5[115]) begin
          axi4Interface_fifoDataBuffer_115 <= s_axis_payload;
        end
        if(_zz_5[116]) begin
          axi4Interface_fifoDataBuffer_116 <= s_axis_payload;
        end
        if(_zz_5[117]) begin
          axi4Interface_fifoDataBuffer_117 <= s_axis_payload;
        end
        if(_zz_5[118]) begin
          axi4Interface_fifoDataBuffer_118 <= s_axis_payload;
        end
        if(_zz_5[119]) begin
          axi4Interface_fifoDataBuffer_119 <= s_axis_payload;
        end
        if(_zz_5[120]) begin
          axi4Interface_fifoDataBuffer_120 <= s_axis_payload;
        end
        if(_zz_5[121]) begin
          axi4Interface_fifoDataBuffer_121 <= s_axis_payload;
        end
        if(_zz_5[122]) begin
          axi4Interface_fifoDataBuffer_122 <= s_axis_payload;
        end
        if(_zz_5[123]) begin
          axi4Interface_fifoDataBuffer_123 <= s_axis_payload;
        end
        if(_zz_5[124]) begin
          axi4Interface_fifoDataBuffer_124 <= s_axis_payload;
        end
        if(_zz_5[125]) begin
          axi4Interface_fifoDataBuffer_125 <= s_axis_payload;
        end
        if(_zz_5[126]) begin
          axi4Interface_fifoDataBuffer_126 <= s_axis_payload;
        end
        if(_zz_5[127]) begin
          axi4Interface_fifoDataBuffer_127 <= s_axis_payload;
        end
        if(_zz_5[128]) begin
          axi4Interface_fifoDataBuffer_128 <= s_axis_payload;
        end
        if(_zz_5[129]) begin
          axi4Interface_fifoDataBuffer_129 <= s_axis_payload;
        end
        if(_zz_5[130]) begin
          axi4Interface_fifoDataBuffer_130 <= s_axis_payload;
        end
        if(_zz_5[131]) begin
          axi4Interface_fifoDataBuffer_131 <= s_axis_payload;
        end
        if(_zz_5[132]) begin
          axi4Interface_fifoDataBuffer_132 <= s_axis_payload;
        end
        if(_zz_5[133]) begin
          axi4Interface_fifoDataBuffer_133 <= s_axis_payload;
        end
        if(_zz_5[134]) begin
          axi4Interface_fifoDataBuffer_134 <= s_axis_payload;
        end
        if(_zz_5[135]) begin
          axi4Interface_fifoDataBuffer_135 <= s_axis_payload;
        end
        if(_zz_5[136]) begin
          axi4Interface_fifoDataBuffer_136 <= s_axis_payload;
        end
        if(_zz_5[137]) begin
          axi4Interface_fifoDataBuffer_137 <= s_axis_payload;
        end
        if(_zz_5[138]) begin
          axi4Interface_fifoDataBuffer_138 <= s_axis_payload;
        end
        if(_zz_5[139]) begin
          axi4Interface_fifoDataBuffer_139 <= s_axis_payload;
        end
        if(_zz_5[140]) begin
          axi4Interface_fifoDataBuffer_140 <= s_axis_payload;
        end
        if(_zz_5[141]) begin
          axi4Interface_fifoDataBuffer_141 <= s_axis_payload;
        end
        if(_zz_5[142]) begin
          axi4Interface_fifoDataBuffer_142 <= s_axis_payload;
        end
        if(_zz_5[143]) begin
          axi4Interface_fifoDataBuffer_143 <= s_axis_payload;
        end
        if(_zz_5[144]) begin
          axi4Interface_fifoDataBuffer_144 <= s_axis_payload;
        end
        if(_zz_5[145]) begin
          axi4Interface_fifoDataBuffer_145 <= s_axis_payload;
        end
        if(_zz_5[146]) begin
          axi4Interface_fifoDataBuffer_146 <= s_axis_payload;
        end
        if(_zz_5[147]) begin
          axi4Interface_fifoDataBuffer_147 <= s_axis_payload;
        end
        if(_zz_5[148]) begin
          axi4Interface_fifoDataBuffer_148 <= s_axis_payload;
        end
        if(_zz_5[149]) begin
          axi4Interface_fifoDataBuffer_149 <= s_axis_payload;
        end
        if(_zz_5[150]) begin
          axi4Interface_fifoDataBuffer_150 <= s_axis_payload;
        end
        if(_zz_5[151]) begin
          axi4Interface_fifoDataBuffer_151 <= s_axis_payload;
        end
        if(_zz_5[152]) begin
          axi4Interface_fifoDataBuffer_152 <= s_axis_payload;
        end
        if(_zz_5[153]) begin
          axi4Interface_fifoDataBuffer_153 <= s_axis_payload;
        end
        if(_zz_5[154]) begin
          axi4Interface_fifoDataBuffer_154 <= s_axis_payload;
        end
        if(_zz_5[155]) begin
          axi4Interface_fifoDataBuffer_155 <= s_axis_payload;
        end
        if(_zz_5[156]) begin
          axi4Interface_fifoDataBuffer_156 <= s_axis_payload;
        end
        if(_zz_5[157]) begin
          axi4Interface_fifoDataBuffer_157 <= s_axis_payload;
        end
        if(_zz_5[158]) begin
          axi4Interface_fifoDataBuffer_158 <= s_axis_payload;
        end
        if(_zz_5[159]) begin
          axi4Interface_fifoDataBuffer_159 <= s_axis_payload;
        end
        if(_zz_5[160]) begin
          axi4Interface_fifoDataBuffer_160 <= s_axis_payload;
        end
        if(_zz_5[161]) begin
          axi4Interface_fifoDataBuffer_161 <= s_axis_payload;
        end
        if(_zz_5[162]) begin
          axi4Interface_fifoDataBuffer_162 <= s_axis_payload;
        end
        if(_zz_5[163]) begin
          axi4Interface_fifoDataBuffer_163 <= s_axis_payload;
        end
        if(_zz_5[164]) begin
          axi4Interface_fifoDataBuffer_164 <= s_axis_payload;
        end
        if(_zz_5[165]) begin
          axi4Interface_fifoDataBuffer_165 <= s_axis_payload;
        end
        if(_zz_5[166]) begin
          axi4Interface_fifoDataBuffer_166 <= s_axis_payload;
        end
        if(_zz_5[167]) begin
          axi4Interface_fifoDataBuffer_167 <= s_axis_payload;
        end
        if(_zz_5[168]) begin
          axi4Interface_fifoDataBuffer_168 <= s_axis_payload;
        end
        if(_zz_5[169]) begin
          axi4Interface_fifoDataBuffer_169 <= s_axis_payload;
        end
        if(_zz_5[170]) begin
          axi4Interface_fifoDataBuffer_170 <= s_axis_payload;
        end
        if(_zz_5[171]) begin
          axi4Interface_fifoDataBuffer_171 <= s_axis_payload;
        end
        if(_zz_5[172]) begin
          axi4Interface_fifoDataBuffer_172 <= s_axis_payload;
        end
        if(_zz_5[173]) begin
          axi4Interface_fifoDataBuffer_173 <= s_axis_payload;
        end
        if(_zz_5[174]) begin
          axi4Interface_fifoDataBuffer_174 <= s_axis_payload;
        end
        if(_zz_5[175]) begin
          axi4Interface_fifoDataBuffer_175 <= s_axis_payload;
        end
        if(_zz_5[176]) begin
          axi4Interface_fifoDataBuffer_176 <= s_axis_payload;
        end
        if(_zz_5[177]) begin
          axi4Interface_fifoDataBuffer_177 <= s_axis_payload;
        end
        if(_zz_5[178]) begin
          axi4Interface_fifoDataBuffer_178 <= s_axis_payload;
        end
        if(_zz_5[179]) begin
          axi4Interface_fifoDataBuffer_179 <= s_axis_payload;
        end
        if(_zz_5[180]) begin
          axi4Interface_fifoDataBuffer_180 <= s_axis_payload;
        end
        if(_zz_5[181]) begin
          axi4Interface_fifoDataBuffer_181 <= s_axis_payload;
        end
        if(_zz_5[182]) begin
          axi4Interface_fifoDataBuffer_182 <= s_axis_payload;
        end
        if(_zz_5[183]) begin
          axi4Interface_fifoDataBuffer_183 <= s_axis_payload;
        end
        if(_zz_5[184]) begin
          axi4Interface_fifoDataBuffer_184 <= s_axis_payload;
        end
        if(_zz_5[185]) begin
          axi4Interface_fifoDataBuffer_185 <= s_axis_payload;
        end
        if(_zz_5[186]) begin
          axi4Interface_fifoDataBuffer_186 <= s_axis_payload;
        end
        if(_zz_5[187]) begin
          axi4Interface_fifoDataBuffer_187 <= s_axis_payload;
        end
        if(_zz_5[188]) begin
          axi4Interface_fifoDataBuffer_188 <= s_axis_payload;
        end
        if(_zz_5[189]) begin
          axi4Interface_fifoDataBuffer_189 <= s_axis_payload;
        end
        if(_zz_5[190]) begin
          axi4Interface_fifoDataBuffer_190 <= s_axis_payload;
        end
        if(_zz_5[191]) begin
          axi4Interface_fifoDataBuffer_191 <= s_axis_payload;
        end
        if(_zz_5[192]) begin
          axi4Interface_fifoDataBuffer_192 <= s_axis_payload;
        end
        if(_zz_5[193]) begin
          axi4Interface_fifoDataBuffer_193 <= s_axis_payload;
        end
        if(_zz_5[194]) begin
          axi4Interface_fifoDataBuffer_194 <= s_axis_payload;
        end
        if(_zz_5[195]) begin
          axi4Interface_fifoDataBuffer_195 <= s_axis_payload;
        end
        if(_zz_5[196]) begin
          axi4Interface_fifoDataBuffer_196 <= s_axis_payload;
        end
        if(_zz_5[197]) begin
          axi4Interface_fifoDataBuffer_197 <= s_axis_payload;
        end
        if(_zz_5[198]) begin
          axi4Interface_fifoDataBuffer_198 <= s_axis_payload;
        end
        if(_zz_5[199]) begin
          axi4Interface_fifoDataBuffer_199 <= s_axis_payload;
        end
        if(_zz_5[200]) begin
          axi4Interface_fifoDataBuffer_200 <= s_axis_payload;
        end
        if(_zz_5[201]) begin
          axi4Interface_fifoDataBuffer_201 <= s_axis_payload;
        end
        if(_zz_5[202]) begin
          axi4Interface_fifoDataBuffer_202 <= s_axis_payload;
        end
        if(_zz_5[203]) begin
          axi4Interface_fifoDataBuffer_203 <= s_axis_payload;
        end
        if(_zz_5[204]) begin
          axi4Interface_fifoDataBuffer_204 <= s_axis_payload;
        end
        if(_zz_5[205]) begin
          axi4Interface_fifoDataBuffer_205 <= s_axis_payload;
        end
        if(_zz_5[206]) begin
          axi4Interface_fifoDataBuffer_206 <= s_axis_payload;
        end
        if(_zz_5[207]) begin
          axi4Interface_fifoDataBuffer_207 <= s_axis_payload;
        end
        if(_zz_5[208]) begin
          axi4Interface_fifoDataBuffer_208 <= s_axis_payload;
        end
        if(_zz_5[209]) begin
          axi4Interface_fifoDataBuffer_209 <= s_axis_payload;
        end
        if(_zz_5[210]) begin
          axi4Interface_fifoDataBuffer_210 <= s_axis_payload;
        end
        if(_zz_5[211]) begin
          axi4Interface_fifoDataBuffer_211 <= s_axis_payload;
        end
        if(_zz_5[212]) begin
          axi4Interface_fifoDataBuffer_212 <= s_axis_payload;
        end
        if(_zz_5[213]) begin
          axi4Interface_fifoDataBuffer_213 <= s_axis_payload;
        end
        if(_zz_5[214]) begin
          axi4Interface_fifoDataBuffer_214 <= s_axis_payload;
        end
        if(_zz_5[215]) begin
          axi4Interface_fifoDataBuffer_215 <= s_axis_payload;
        end
        if(_zz_5[216]) begin
          axi4Interface_fifoDataBuffer_216 <= s_axis_payload;
        end
        if(_zz_5[217]) begin
          axi4Interface_fifoDataBuffer_217 <= s_axis_payload;
        end
        if(_zz_5[218]) begin
          axi4Interface_fifoDataBuffer_218 <= s_axis_payload;
        end
        if(_zz_5[219]) begin
          axi4Interface_fifoDataBuffer_219 <= s_axis_payload;
        end
        if(_zz_5[220]) begin
          axi4Interface_fifoDataBuffer_220 <= s_axis_payload;
        end
        if(_zz_5[221]) begin
          axi4Interface_fifoDataBuffer_221 <= s_axis_payload;
        end
        if(_zz_5[222]) begin
          axi4Interface_fifoDataBuffer_222 <= s_axis_payload;
        end
        if(_zz_5[223]) begin
          axi4Interface_fifoDataBuffer_223 <= s_axis_payload;
        end
        if(_zz_5[224]) begin
          axi4Interface_fifoDataBuffer_224 <= s_axis_payload;
        end
        if(_zz_5[225]) begin
          axi4Interface_fifoDataBuffer_225 <= s_axis_payload;
        end
        if(_zz_5[226]) begin
          axi4Interface_fifoDataBuffer_226 <= s_axis_payload;
        end
        if(_zz_5[227]) begin
          axi4Interface_fifoDataBuffer_227 <= s_axis_payload;
        end
        if(_zz_5[228]) begin
          axi4Interface_fifoDataBuffer_228 <= s_axis_payload;
        end
        if(_zz_5[229]) begin
          axi4Interface_fifoDataBuffer_229 <= s_axis_payload;
        end
        if(_zz_5[230]) begin
          axi4Interface_fifoDataBuffer_230 <= s_axis_payload;
        end
        if(_zz_5[231]) begin
          axi4Interface_fifoDataBuffer_231 <= s_axis_payload;
        end
        if(_zz_5[232]) begin
          axi4Interface_fifoDataBuffer_232 <= s_axis_payload;
        end
        if(_zz_5[233]) begin
          axi4Interface_fifoDataBuffer_233 <= s_axis_payload;
        end
        if(_zz_5[234]) begin
          axi4Interface_fifoDataBuffer_234 <= s_axis_payload;
        end
        if(_zz_5[235]) begin
          axi4Interface_fifoDataBuffer_235 <= s_axis_payload;
        end
        if(_zz_5[236]) begin
          axi4Interface_fifoDataBuffer_236 <= s_axis_payload;
        end
        if(_zz_5[237]) begin
          axi4Interface_fifoDataBuffer_237 <= s_axis_payload;
        end
        if(_zz_5[238]) begin
          axi4Interface_fifoDataBuffer_238 <= s_axis_payload;
        end
        if(_zz_5[239]) begin
          axi4Interface_fifoDataBuffer_239 <= s_axis_payload;
        end
        if(_zz_5[240]) begin
          axi4Interface_fifoDataBuffer_240 <= s_axis_payload;
        end
        if(_zz_5[241]) begin
          axi4Interface_fifoDataBuffer_241 <= s_axis_payload;
        end
        if(_zz_5[242]) begin
          axi4Interface_fifoDataBuffer_242 <= s_axis_payload;
        end
        if(_zz_5[243]) begin
          axi4Interface_fifoDataBuffer_243 <= s_axis_payload;
        end
        if(_zz_5[244]) begin
          axi4Interface_fifoDataBuffer_244 <= s_axis_payload;
        end
        if(_zz_5[245]) begin
          axi4Interface_fifoDataBuffer_245 <= s_axis_payload;
        end
        if(_zz_5[246]) begin
          axi4Interface_fifoDataBuffer_246 <= s_axis_payload;
        end
        if(_zz_5[247]) begin
          axi4Interface_fifoDataBuffer_247 <= s_axis_payload;
        end
        if(_zz_5[248]) begin
          axi4Interface_fifoDataBuffer_248 <= s_axis_payload;
        end
        if(_zz_5[249]) begin
          axi4Interface_fifoDataBuffer_249 <= s_axis_payload;
        end
        if(_zz_5[250]) begin
          axi4Interface_fifoDataBuffer_250 <= s_axis_payload;
        end
        if(_zz_5[251]) begin
          axi4Interface_fifoDataBuffer_251 <= s_axis_payload;
        end
        if(_zz_5[252]) begin
          axi4Interface_fifoDataBuffer_252 <= s_axis_payload;
        end
        if(_zz_5[253]) begin
          axi4Interface_fifoDataBuffer_253 <= s_axis_payload;
        end
        if(_zz_5[254]) begin
          axi4Interface_fifoDataBuffer_254 <= s_axis_payload;
        end
        if(_zz_5[255]) begin
          axi4Interface_fifoDataBuffer_255 <= s_axis_payload;
        end
      end
      if(axi4Interface_t_w_fire) begin
        axi4Interface_address <= Axi4Incr_result;
      end
      if(aresetn) begin
        axi4Interface_isTransferAfterReset <= 1'b0;
      end
      if(aresetn) begin
        if(axi4Interface_t_aw_fire) begin
          axi4Interface_controlAwValid <= 1'b0;
        end
        if(when_Axi4WriteMaster_l92) begin
          axi4Interface_controlAwValid <= 1'b1;
        end
      end
      if(_zz_when_Axi4WriteMaster_l92) begin
        axi4Interface_initialAddress <= axi4Interface_address;
      end
      if(when_Axi4WriteMaster_l156) begin
        axi4Interface_controlBReady <= 1'b1;
      end
      if(axi4Interface_t_b_fire) begin
        axi4Interface_controlBReady <= 1'b0;
      end
    end
  end

  always @(posedge aclk) begin
    m_axi_wvalid_regNext <= m_axi_wvalid;
  end


endmodule
