// Generator : SpinalHDL v1.5.0    git head : 83a031922866b078c411ec5529e00f1b6e79f8e7
// Component : TestAxi4WriteMaster
// Git hash  : 0979837f915a50e3cecc964d3b3d2423bf347c03



module TestAxi4WriteMaster (
  input               fifoValid,
  output reg          fifoReady,
  input      [31:0]   fifoPayload,
  output              awValid,
  input               awReady,
  output reg [31:0]   awaddr,
  output     [0:0]    awid,
  output     [3:0]    awregion,
  output     [7:0]    awlen,
  output     [2:0]    awsize,
  output     [1:0]    awburst,
  output     [0:0]    awlock,
  output     [3:0]    awcache,
  output     [3:0]    awqos,
  output     [2:0]    awprot,
  output reg          wValid,
  input               wReady,
  output reg [31:0]   wdata,
  output     [3:0]    wstrb,
  output              wlast,
  input               bValid,
  output              bReady,
  input      [0:0]    bid,
  input      [1:0]    bresp,
  output              arValid,
  input               arReady,
  output     [31:0]   araddr,
  output     [0:0]    arid,
  output     [3:0]    arregion,
  output     [7:0]    arlen,
  output     [2:0]    arsize,
  output     [1:0]    arburst,
  output     [0:0]    arlock,
  output     [3:0]    arcache,
  output     [3:0]    arqos,
  output     [2:0]    arprot,
  input               rValid,
  output              rReady,
  input      [31:0]   rdata,
  input      [0:0]    rid,
  input      [1:0]    rresp,
  input               rlast,
  input               clk,
  input               reset
);
  wire       [8:0]    _zz__zz_wdata_1;
  wire       [0:0]    _zz__zz_wdata_1_1;
  wire       [8:0]    _zz__zz_when_Axi4WriteMaster_l53_1;
  wire       [0:0]    _zz__zz_when_Axi4WriteMaster_l53_1_1;
  wire       [7:0]    _zz__zz_5;
  wire       [1:0]    _zz_Axi4Incr_alignMask;
  wire       [11:0]   _zz_Axi4Incr_base;
  wire       [11:0]   _zz_Axi4Incr_base_1;
  wire       [11:0]   _zz_Axi4Incr_baseIncr;
  wire       [2:0]    _zz_Axi4Incr_wrapCase_1;
  wire       [2:0]    _zz_Axi4Incr_wrapCase_2;
  reg        [11:0]   _zz_Axi4Incr_result;
  wire       [10:0]   _zz_Axi4Incr_result_1;
  wire       [0:0]    _zz_Axi4Incr_result_2;
  wire       [9:0]    _zz_Axi4Incr_result_3;
  wire       [1:0]    _zz_Axi4Incr_result_4;
  wire       [8:0]    _zz_Axi4Incr_result_5;
  wire       [2:0]    _zz_Axi4Incr_result_6;
  wire       [7:0]    _zz_Axi4Incr_result_7;
  wire       [3:0]    _zz_Axi4Incr_result_8;
  wire       [6:0]    _zz_Axi4Incr_result_9;
  wire       [4:0]    _zz_Axi4Incr_result_10;
  wire       [5:0]    _zz_Axi4Incr_result_11;
  wire       [5:0]    _zz_Axi4Incr_result_12;
  reg        [31:0]   _zz_wdata_3;
  wire       [7:0]    _zz_wdata_4;
  reg                 _zz_wdata;
  reg                 _zz_1;
  reg        [8:0]    _zz_wdata_1;
  reg        [8:0]    _zz_wdata_2;
  wire                _zz_when_Axi4WriteMaster_l61;
  wire                _zz_2;
  reg                 _zz_when_Axi4WriteMaster_l53;
  reg                 _zz_3;
  reg        [8:0]    _zz_when_Axi4WriteMaster_l53_1;
  reg        [8:0]    _zz_when_Axi4WriteMaster_l53_2;
  wire                _zz_when_Axi4WriteMaster_l53_3;
  wire                _zz_4;
  reg        [31:0]   fifoDataBuffer_0;
  reg        [31:0]   fifoDataBuffer_1;
  reg        [31:0]   fifoDataBuffer_2;
  reg        [31:0]   fifoDataBuffer_3;
  reg        [31:0]   fifoDataBuffer_4;
  reg        [31:0]   fifoDataBuffer_5;
  reg        [31:0]   fifoDataBuffer_6;
  reg        [31:0]   fifoDataBuffer_7;
  reg        [31:0]   fifoDataBuffer_8;
  reg        [31:0]   fifoDataBuffer_9;
  reg        [31:0]   fifoDataBuffer_10;
  reg        [31:0]   fifoDataBuffer_11;
  reg        [31:0]   fifoDataBuffer_12;
  reg        [31:0]   fifoDataBuffer_13;
  reg        [31:0]   fifoDataBuffer_14;
  reg        [31:0]   fifoDataBuffer_15;
  reg        [31:0]   fifoDataBuffer_16;
  reg        [31:0]   fifoDataBuffer_17;
  reg        [31:0]   fifoDataBuffer_18;
  reg        [31:0]   fifoDataBuffer_19;
  reg        [31:0]   fifoDataBuffer_20;
  reg        [31:0]   fifoDataBuffer_21;
  reg        [31:0]   fifoDataBuffer_22;
  reg        [31:0]   fifoDataBuffer_23;
  reg        [31:0]   fifoDataBuffer_24;
  reg        [31:0]   fifoDataBuffer_25;
  reg        [31:0]   fifoDataBuffer_26;
  reg        [31:0]   fifoDataBuffer_27;
  reg        [31:0]   fifoDataBuffer_28;
  reg        [31:0]   fifoDataBuffer_29;
  reg        [31:0]   fifoDataBuffer_30;
  reg        [31:0]   fifoDataBuffer_31;
  reg        [31:0]   fifoDataBuffer_32;
  reg        [31:0]   fifoDataBuffer_33;
  reg        [31:0]   fifoDataBuffer_34;
  reg        [31:0]   fifoDataBuffer_35;
  reg        [31:0]   fifoDataBuffer_36;
  reg        [31:0]   fifoDataBuffer_37;
  reg        [31:0]   fifoDataBuffer_38;
  reg        [31:0]   fifoDataBuffer_39;
  reg        [31:0]   fifoDataBuffer_40;
  reg        [31:0]   fifoDataBuffer_41;
  reg        [31:0]   fifoDataBuffer_42;
  reg        [31:0]   fifoDataBuffer_43;
  reg        [31:0]   fifoDataBuffer_44;
  reg        [31:0]   fifoDataBuffer_45;
  reg        [31:0]   fifoDataBuffer_46;
  reg        [31:0]   fifoDataBuffer_47;
  reg        [31:0]   fifoDataBuffer_48;
  reg        [31:0]   fifoDataBuffer_49;
  reg        [31:0]   fifoDataBuffer_50;
  reg        [31:0]   fifoDataBuffer_51;
  reg        [31:0]   fifoDataBuffer_52;
  reg        [31:0]   fifoDataBuffer_53;
  reg        [31:0]   fifoDataBuffer_54;
  reg        [31:0]   fifoDataBuffer_55;
  reg        [31:0]   fifoDataBuffer_56;
  reg        [31:0]   fifoDataBuffer_57;
  reg        [31:0]   fifoDataBuffer_58;
  reg        [31:0]   fifoDataBuffer_59;
  reg        [31:0]   fifoDataBuffer_60;
  reg        [31:0]   fifoDataBuffer_61;
  reg        [31:0]   fifoDataBuffer_62;
  reg        [31:0]   fifoDataBuffer_63;
  reg        [31:0]   fifoDataBuffer_64;
  reg        [31:0]   fifoDataBuffer_65;
  reg        [31:0]   fifoDataBuffer_66;
  reg        [31:0]   fifoDataBuffer_67;
  reg        [31:0]   fifoDataBuffer_68;
  reg        [31:0]   fifoDataBuffer_69;
  reg        [31:0]   fifoDataBuffer_70;
  reg        [31:0]   fifoDataBuffer_71;
  reg        [31:0]   fifoDataBuffer_72;
  reg        [31:0]   fifoDataBuffer_73;
  reg        [31:0]   fifoDataBuffer_74;
  reg        [31:0]   fifoDataBuffer_75;
  reg        [31:0]   fifoDataBuffer_76;
  reg        [31:0]   fifoDataBuffer_77;
  reg        [31:0]   fifoDataBuffer_78;
  reg        [31:0]   fifoDataBuffer_79;
  reg        [31:0]   fifoDataBuffer_80;
  reg        [31:0]   fifoDataBuffer_81;
  reg        [31:0]   fifoDataBuffer_82;
  reg        [31:0]   fifoDataBuffer_83;
  reg        [31:0]   fifoDataBuffer_84;
  reg        [31:0]   fifoDataBuffer_85;
  reg        [31:0]   fifoDataBuffer_86;
  reg        [31:0]   fifoDataBuffer_87;
  reg        [31:0]   fifoDataBuffer_88;
  reg        [31:0]   fifoDataBuffer_89;
  reg        [31:0]   fifoDataBuffer_90;
  reg        [31:0]   fifoDataBuffer_91;
  reg        [31:0]   fifoDataBuffer_92;
  reg        [31:0]   fifoDataBuffer_93;
  reg        [31:0]   fifoDataBuffer_94;
  reg        [31:0]   fifoDataBuffer_95;
  reg        [31:0]   fifoDataBuffer_96;
  reg        [31:0]   fifoDataBuffer_97;
  reg        [31:0]   fifoDataBuffer_98;
  reg        [31:0]   fifoDataBuffer_99;
  reg        [31:0]   fifoDataBuffer_100;
  reg        [31:0]   fifoDataBuffer_101;
  reg        [31:0]   fifoDataBuffer_102;
  reg        [31:0]   fifoDataBuffer_103;
  reg        [31:0]   fifoDataBuffer_104;
  reg        [31:0]   fifoDataBuffer_105;
  reg        [31:0]   fifoDataBuffer_106;
  reg        [31:0]   fifoDataBuffer_107;
  reg        [31:0]   fifoDataBuffer_108;
  reg        [31:0]   fifoDataBuffer_109;
  reg        [31:0]   fifoDataBuffer_110;
  reg        [31:0]   fifoDataBuffer_111;
  reg        [31:0]   fifoDataBuffer_112;
  reg        [31:0]   fifoDataBuffer_113;
  reg        [31:0]   fifoDataBuffer_114;
  reg        [31:0]   fifoDataBuffer_115;
  reg        [31:0]   fifoDataBuffer_116;
  reg        [31:0]   fifoDataBuffer_117;
  reg        [31:0]   fifoDataBuffer_118;
  reg        [31:0]   fifoDataBuffer_119;
  reg        [31:0]   fifoDataBuffer_120;
  reg        [31:0]   fifoDataBuffer_121;
  reg        [31:0]   fifoDataBuffer_122;
  reg        [31:0]   fifoDataBuffer_123;
  reg        [31:0]   fifoDataBuffer_124;
  reg        [31:0]   fifoDataBuffer_125;
  reg        [31:0]   fifoDataBuffer_126;
  reg        [31:0]   fifoDataBuffer_127;
  reg        [31:0]   fifoDataBuffer_128;
  reg        [31:0]   fifoDataBuffer_129;
  reg        [31:0]   fifoDataBuffer_130;
  reg        [31:0]   fifoDataBuffer_131;
  reg        [31:0]   fifoDataBuffer_132;
  reg        [31:0]   fifoDataBuffer_133;
  reg        [31:0]   fifoDataBuffer_134;
  reg        [31:0]   fifoDataBuffer_135;
  reg        [31:0]   fifoDataBuffer_136;
  reg        [31:0]   fifoDataBuffer_137;
  reg        [31:0]   fifoDataBuffer_138;
  reg        [31:0]   fifoDataBuffer_139;
  reg        [31:0]   fifoDataBuffer_140;
  reg        [31:0]   fifoDataBuffer_141;
  reg        [31:0]   fifoDataBuffer_142;
  reg        [31:0]   fifoDataBuffer_143;
  reg        [31:0]   fifoDataBuffer_144;
  reg        [31:0]   fifoDataBuffer_145;
  reg        [31:0]   fifoDataBuffer_146;
  reg        [31:0]   fifoDataBuffer_147;
  reg        [31:0]   fifoDataBuffer_148;
  reg        [31:0]   fifoDataBuffer_149;
  reg        [31:0]   fifoDataBuffer_150;
  reg        [31:0]   fifoDataBuffer_151;
  reg        [31:0]   fifoDataBuffer_152;
  reg        [31:0]   fifoDataBuffer_153;
  reg        [31:0]   fifoDataBuffer_154;
  reg        [31:0]   fifoDataBuffer_155;
  reg        [31:0]   fifoDataBuffer_156;
  reg        [31:0]   fifoDataBuffer_157;
  reg        [31:0]   fifoDataBuffer_158;
  reg        [31:0]   fifoDataBuffer_159;
  reg        [31:0]   fifoDataBuffer_160;
  reg        [31:0]   fifoDataBuffer_161;
  reg        [31:0]   fifoDataBuffer_162;
  reg        [31:0]   fifoDataBuffer_163;
  reg        [31:0]   fifoDataBuffer_164;
  reg        [31:0]   fifoDataBuffer_165;
  reg        [31:0]   fifoDataBuffer_166;
  reg        [31:0]   fifoDataBuffer_167;
  reg        [31:0]   fifoDataBuffer_168;
  reg        [31:0]   fifoDataBuffer_169;
  reg        [31:0]   fifoDataBuffer_170;
  reg        [31:0]   fifoDataBuffer_171;
  reg        [31:0]   fifoDataBuffer_172;
  reg        [31:0]   fifoDataBuffer_173;
  reg        [31:0]   fifoDataBuffer_174;
  reg        [31:0]   fifoDataBuffer_175;
  reg        [31:0]   fifoDataBuffer_176;
  reg        [31:0]   fifoDataBuffer_177;
  reg        [31:0]   fifoDataBuffer_178;
  reg        [31:0]   fifoDataBuffer_179;
  reg        [31:0]   fifoDataBuffer_180;
  reg        [31:0]   fifoDataBuffer_181;
  reg        [31:0]   fifoDataBuffer_182;
  reg        [31:0]   fifoDataBuffer_183;
  reg        [31:0]   fifoDataBuffer_184;
  reg        [31:0]   fifoDataBuffer_185;
  reg        [31:0]   fifoDataBuffer_186;
  reg        [31:0]   fifoDataBuffer_187;
  reg        [31:0]   fifoDataBuffer_188;
  reg        [31:0]   fifoDataBuffer_189;
  reg        [31:0]   fifoDataBuffer_190;
  reg        [31:0]   fifoDataBuffer_191;
  reg        [31:0]   fifoDataBuffer_192;
  reg        [31:0]   fifoDataBuffer_193;
  reg        [31:0]   fifoDataBuffer_194;
  reg        [31:0]   fifoDataBuffer_195;
  reg        [31:0]   fifoDataBuffer_196;
  reg        [31:0]   fifoDataBuffer_197;
  reg        [31:0]   fifoDataBuffer_198;
  reg        [31:0]   fifoDataBuffer_199;
  reg        [31:0]   fifoDataBuffer_200;
  reg        [31:0]   fifoDataBuffer_201;
  reg        [31:0]   fifoDataBuffer_202;
  reg        [31:0]   fifoDataBuffer_203;
  reg        [31:0]   fifoDataBuffer_204;
  reg        [31:0]   fifoDataBuffer_205;
  reg        [31:0]   fifoDataBuffer_206;
  reg        [31:0]   fifoDataBuffer_207;
  reg        [31:0]   fifoDataBuffer_208;
  reg        [31:0]   fifoDataBuffer_209;
  reg        [31:0]   fifoDataBuffer_210;
  reg        [31:0]   fifoDataBuffer_211;
  reg        [31:0]   fifoDataBuffer_212;
  reg        [31:0]   fifoDataBuffer_213;
  reg        [31:0]   fifoDataBuffer_214;
  reg        [31:0]   fifoDataBuffer_215;
  reg        [31:0]   fifoDataBuffer_216;
  reg        [31:0]   fifoDataBuffer_217;
  reg        [31:0]   fifoDataBuffer_218;
  reg        [31:0]   fifoDataBuffer_219;
  reg        [31:0]   fifoDataBuffer_220;
  reg        [31:0]   fifoDataBuffer_221;
  reg        [31:0]   fifoDataBuffer_222;
  reg        [31:0]   fifoDataBuffer_223;
  reg        [31:0]   fifoDataBuffer_224;
  reg        [31:0]   fifoDataBuffer_225;
  reg        [31:0]   fifoDataBuffer_226;
  reg        [31:0]   fifoDataBuffer_227;
  reg        [31:0]   fifoDataBuffer_228;
  reg        [31:0]   fifoDataBuffer_229;
  reg        [31:0]   fifoDataBuffer_230;
  reg        [31:0]   fifoDataBuffer_231;
  reg        [31:0]   fifoDataBuffer_232;
  reg        [31:0]   fifoDataBuffer_233;
  reg        [31:0]   fifoDataBuffer_234;
  reg        [31:0]   fifoDataBuffer_235;
  reg        [31:0]   fifoDataBuffer_236;
  reg        [31:0]   fifoDataBuffer_237;
  reg        [31:0]   fifoDataBuffer_238;
  reg        [31:0]   fifoDataBuffer_239;
  reg        [31:0]   fifoDataBuffer_240;
  reg        [31:0]   fifoDataBuffer_241;
  reg        [31:0]   fifoDataBuffer_242;
  reg        [31:0]   fifoDataBuffer_243;
  reg        [31:0]   fifoDataBuffer_244;
  reg        [31:0]   fifoDataBuffer_245;
  reg        [31:0]   fifoDataBuffer_246;
  reg        [31:0]   fifoDataBuffer_247;
  reg        [31:0]   fifoDataBuffer_248;
  reg        [31:0]   fifoDataBuffer_249;
  reg        [31:0]   fifoDataBuffer_250;
  reg        [31:0]   fifoDataBuffer_251;
  reg        [31:0]   fifoDataBuffer_252;
  reg        [31:0]   fifoDataBuffer_253;
  reg        [31:0]   fifoDataBuffer_254;
  reg        [31:0]   fifoDataBuffer_255;
  wire                when_Axi4WriteMaster_l47;
  wire       [255:0]  _zz_5;
  wire                when_Axi4WriteMaster_l53;
  wire                when_Axi4WriteMaster_l61;
  reg        [31:0]   axi4Interface_address;
  wire                when_Axi4WriteMaster_l70;
  wire       [1:0]    Axi4Incr_validSize;
  reg        [31:0]   Axi4Incr_result;
  wire       [19:0]   Axi4Incr_highCat;
  wire       [2:0]    Axi4Incr_sizeValue;
  wire       [11:0]   Axi4Incr_alignMask;
  wire       [11:0]   Axi4Incr_base;
  wire       [11:0]   Axi4Incr_baseIncr;
  reg        [1:0]    _zz_Axi4Incr_wrapCase;
  wire       [2:0]    Axi4Incr_wrapCase;
  reg        [31:0]   axi4Interface_initialAddress;
  wire                when_Axi4WriteMaster_l87;
  wire                when_Axi4WriteMaster_l118;
  wire                when_Axi4WriteMaster_l124;

  assign _zz__zz_wdata_1_1 = _zz_wdata;
  assign _zz__zz_wdata_1 = {8'd0, _zz__zz_wdata_1_1};
  assign _zz__zz_when_Axi4WriteMaster_l53_1_1 = _zz_when_Axi4WriteMaster_l53;
  assign _zz__zz_when_Axi4WriteMaster_l53_1 = {8'd0, _zz__zz_when_Axi4WriteMaster_l53_1_1};
  assign _zz__zz_5 = _zz_when_Axi4WriteMaster_l53_2[7:0];
  assign _zz_Axi4Incr_alignMask = {(2'b01 < Axi4Incr_validSize),(2'b00 < Axi4Incr_validSize)};
  assign _zz_Axi4Incr_base_1 = axi4Interface_address[11 : 0];
  assign _zz_Axi4Incr_base = _zz_Axi4Incr_base_1;
  assign _zz_Axi4Incr_baseIncr = {9'd0, Axi4Incr_sizeValue};
  assign _zz_Axi4Incr_wrapCase_1 = {1'd0, Axi4Incr_validSize};
  assign _zz_Axi4Incr_wrapCase_2 = {1'd0, _zz_Axi4Incr_wrapCase};
  assign _zz_wdata_4 = _zz_wdata_2[7:0];
  assign _zz_Axi4Incr_result_1 = Axi4Incr_base[11 : 1];
  assign _zz_Axi4Incr_result_2 = Axi4Incr_baseIncr[0 : 0];
  assign _zz_Axi4Incr_result_3 = Axi4Incr_base[11 : 2];
  assign _zz_Axi4Incr_result_4 = Axi4Incr_baseIncr[1 : 0];
  assign _zz_Axi4Incr_result_5 = Axi4Incr_base[11 : 3];
  assign _zz_Axi4Incr_result_6 = Axi4Incr_baseIncr[2 : 0];
  assign _zz_Axi4Incr_result_7 = Axi4Incr_base[11 : 4];
  assign _zz_Axi4Incr_result_8 = Axi4Incr_baseIncr[3 : 0];
  assign _zz_Axi4Incr_result_9 = Axi4Incr_base[11 : 5];
  assign _zz_Axi4Incr_result_10 = Axi4Incr_baseIncr[4 : 0];
  assign _zz_Axi4Incr_result_11 = Axi4Incr_base[11 : 6];
  assign _zz_Axi4Incr_result_12 = Axi4Incr_baseIncr[5 : 0];
  always @(*) begin
    case(Axi4Incr_wrapCase)
      3'b000 : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_1,_zz_Axi4Incr_result_2};
      end
      3'b001 : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_3,_zz_Axi4Incr_result_4};
      end
      3'b010 : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_5,_zz_Axi4Incr_result_6};
      end
      3'b011 : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_7,_zz_Axi4Incr_result_8};
      end
      3'b100 : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_9,_zz_Axi4Incr_result_10};
      end
      default : begin
        _zz_Axi4Incr_result = {_zz_Axi4Incr_result_11,_zz_Axi4Incr_result_12};
      end
    endcase
  end

  always @(*) begin
    case(_zz_wdata_4)
      8'b00000000 : begin
        _zz_wdata_3 = fifoDataBuffer_0;
      end
      8'b00000001 : begin
        _zz_wdata_3 = fifoDataBuffer_1;
      end
      8'b00000010 : begin
        _zz_wdata_3 = fifoDataBuffer_2;
      end
      8'b00000011 : begin
        _zz_wdata_3 = fifoDataBuffer_3;
      end
      8'b00000100 : begin
        _zz_wdata_3 = fifoDataBuffer_4;
      end
      8'b00000101 : begin
        _zz_wdata_3 = fifoDataBuffer_5;
      end
      8'b00000110 : begin
        _zz_wdata_3 = fifoDataBuffer_6;
      end
      8'b00000111 : begin
        _zz_wdata_3 = fifoDataBuffer_7;
      end
      8'b00001000 : begin
        _zz_wdata_3 = fifoDataBuffer_8;
      end
      8'b00001001 : begin
        _zz_wdata_3 = fifoDataBuffer_9;
      end
      8'b00001010 : begin
        _zz_wdata_3 = fifoDataBuffer_10;
      end
      8'b00001011 : begin
        _zz_wdata_3 = fifoDataBuffer_11;
      end
      8'b00001100 : begin
        _zz_wdata_3 = fifoDataBuffer_12;
      end
      8'b00001101 : begin
        _zz_wdata_3 = fifoDataBuffer_13;
      end
      8'b00001110 : begin
        _zz_wdata_3 = fifoDataBuffer_14;
      end
      8'b00001111 : begin
        _zz_wdata_3 = fifoDataBuffer_15;
      end
      8'b00010000 : begin
        _zz_wdata_3 = fifoDataBuffer_16;
      end
      8'b00010001 : begin
        _zz_wdata_3 = fifoDataBuffer_17;
      end
      8'b00010010 : begin
        _zz_wdata_3 = fifoDataBuffer_18;
      end
      8'b00010011 : begin
        _zz_wdata_3 = fifoDataBuffer_19;
      end
      8'b00010100 : begin
        _zz_wdata_3 = fifoDataBuffer_20;
      end
      8'b00010101 : begin
        _zz_wdata_3 = fifoDataBuffer_21;
      end
      8'b00010110 : begin
        _zz_wdata_3 = fifoDataBuffer_22;
      end
      8'b00010111 : begin
        _zz_wdata_3 = fifoDataBuffer_23;
      end
      8'b00011000 : begin
        _zz_wdata_3 = fifoDataBuffer_24;
      end
      8'b00011001 : begin
        _zz_wdata_3 = fifoDataBuffer_25;
      end
      8'b00011010 : begin
        _zz_wdata_3 = fifoDataBuffer_26;
      end
      8'b00011011 : begin
        _zz_wdata_3 = fifoDataBuffer_27;
      end
      8'b00011100 : begin
        _zz_wdata_3 = fifoDataBuffer_28;
      end
      8'b00011101 : begin
        _zz_wdata_3 = fifoDataBuffer_29;
      end
      8'b00011110 : begin
        _zz_wdata_3 = fifoDataBuffer_30;
      end
      8'b00011111 : begin
        _zz_wdata_3 = fifoDataBuffer_31;
      end
      8'b00100000 : begin
        _zz_wdata_3 = fifoDataBuffer_32;
      end
      8'b00100001 : begin
        _zz_wdata_3 = fifoDataBuffer_33;
      end
      8'b00100010 : begin
        _zz_wdata_3 = fifoDataBuffer_34;
      end
      8'b00100011 : begin
        _zz_wdata_3 = fifoDataBuffer_35;
      end
      8'b00100100 : begin
        _zz_wdata_3 = fifoDataBuffer_36;
      end
      8'b00100101 : begin
        _zz_wdata_3 = fifoDataBuffer_37;
      end
      8'b00100110 : begin
        _zz_wdata_3 = fifoDataBuffer_38;
      end
      8'b00100111 : begin
        _zz_wdata_3 = fifoDataBuffer_39;
      end
      8'b00101000 : begin
        _zz_wdata_3 = fifoDataBuffer_40;
      end
      8'b00101001 : begin
        _zz_wdata_3 = fifoDataBuffer_41;
      end
      8'b00101010 : begin
        _zz_wdata_3 = fifoDataBuffer_42;
      end
      8'b00101011 : begin
        _zz_wdata_3 = fifoDataBuffer_43;
      end
      8'b00101100 : begin
        _zz_wdata_3 = fifoDataBuffer_44;
      end
      8'b00101101 : begin
        _zz_wdata_3 = fifoDataBuffer_45;
      end
      8'b00101110 : begin
        _zz_wdata_3 = fifoDataBuffer_46;
      end
      8'b00101111 : begin
        _zz_wdata_3 = fifoDataBuffer_47;
      end
      8'b00110000 : begin
        _zz_wdata_3 = fifoDataBuffer_48;
      end
      8'b00110001 : begin
        _zz_wdata_3 = fifoDataBuffer_49;
      end
      8'b00110010 : begin
        _zz_wdata_3 = fifoDataBuffer_50;
      end
      8'b00110011 : begin
        _zz_wdata_3 = fifoDataBuffer_51;
      end
      8'b00110100 : begin
        _zz_wdata_3 = fifoDataBuffer_52;
      end
      8'b00110101 : begin
        _zz_wdata_3 = fifoDataBuffer_53;
      end
      8'b00110110 : begin
        _zz_wdata_3 = fifoDataBuffer_54;
      end
      8'b00110111 : begin
        _zz_wdata_3 = fifoDataBuffer_55;
      end
      8'b00111000 : begin
        _zz_wdata_3 = fifoDataBuffer_56;
      end
      8'b00111001 : begin
        _zz_wdata_3 = fifoDataBuffer_57;
      end
      8'b00111010 : begin
        _zz_wdata_3 = fifoDataBuffer_58;
      end
      8'b00111011 : begin
        _zz_wdata_3 = fifoDataBuffer_59;
      end
      8'b00111100 : begin
        _zz_wdata_3 = fifoDataBuffer_60;
      end
      8'b00111101 : begin
        _zz_wdata_3 = fifoDataBuffer_61;
      end
      8'b00111110 : begin
        _zz_wdata_3 = fifoDataBuffer_62;
      end
      8'b00111111 : begin
        _zz_wdata_3 = fifoDataBuffer_63;
      end
      8'b01000000 : begin
        _zz_wdata_3 = fifoDataBuffer_64;
      end
      8'b01000001 : begin
        _zz_wdata_3 = fifoDataBuffer_65;
      end
      8'b01000010 : begin
        _zz_wdata_3 = fifoDataBuffer_66;
      end
      8'b01000011 : begin
        _zz_wdata_3 = fifoDataBuffer_67;
      end
      8'b01000100 : begin
        _zz_wdata_3 = fifoDataBuffer_68;
      end
      8'b01000101 : begin
        _zz_wdata_3 = fifoDataBuffer_69;
      end
      8'b01000110 : begin
        _zz_wdata_3 = fifoDataBuffer_70;
      end
      8'b01000111 : begin
        _zz_wdata_3 = fifoDataBuffer_71;
      end
      8'b01001000 : begin
        _zz_wdata_3 = fifoDataBuffer_72;
      end
      8'b01001001 : begin
        _zz_wdata_3 = fifoDataBuffer_73;
      end
      8'b01001010 : begin
        _zz_wdata_3 = fifoDataBuffer_74;
      end
      8'b01001011 : begin
        _zz_wdata_3 = fifoDataBuffer_75;
      end
      8'b01001100 : begin
        _zz_wdata_3 = fifoDataBuffer_76;
      end
      8'b01001101 : begin
        _zz_wdata_3 = fifoDataBuffer_77;
      end
      8'b01001110 : begin
        _zz_wdata_3 = fifoDataBuffer_78;
      end
      8'b01001111 : begin
        _zz_wdata_3 = fifoDataBuffer_79;
      end
      8'b01010000 : begin
        _zz_wdata_3 = fifoDataBuffer_80;
      end
      8'b01010001 : begin
        _zz_wdata_3 = fifoDataBuffer_81;
      end
      8'b01010010 : begin
        _zz_wdata_3 = fifoDataBuffer_82;
      end
      8'b01010011 : begin
        _zz_wdata_3 = fifoDataBuffer_83;
      end
      8'b01010100 : begin
        _zz_wdata_3 = fifoDataBuffer_84;
      end
      8'b01010101 : begin
        _zz_wdata_3 = fifoDataBuffer_85;
      end
      8'b01010110 : begin
        _zz_wdata_3 = fifoDataBuffer_86;
      end
      8'b01010111 : begin
        _zz_wdata_3 = fifoDataBuffer_87;
      end
      8'b01011000 : begin
        _zz_wdata_3 = fifoDataBuffer_88;
      end
      8'b01011001 : begin
        _zz_wdata_3 = fifoDataBuffer_89;
      end
      8'b01011010 : begin
        _zz_wdata_3 = fifoDataBuffer_90;
      end
      8'b01011011 : begin
        _zz_wdata_3 = fifoDataBuffer_91;
      end
      8'b01011100 : begin
        _zz_wdata_3 = fifoDataBuffer_92;
      end
      8'b01011101 : begin
        _zz_wdata_3 = fifoDataBuffer_93;
      end
      8'b01011110 : begin
        _zz_wdata_3 = fifoDataBuffer_94;
      end
      8'b01011111 : begin
        _zz_wdata_3 = fifoDataBuffer_95;
      end
      8'b01100000 : begin
        _zz_wdata_3 = fifoDataBuffer_96;
      end
      8'b01100001 : begin
        _zz_wdata_3 = fifoDataBuffer_97;
      end
      8'b01100010 : begin
        _zz_wdata_3 = fifoDataBuffer_98;
      end
      8'b01100011 : begin
        _zz_wdata_3 = fifoDataBuffer_99;
      end
      8'b01100100 : begin
        _zz_wdata_3 = fifoDataBuffer_100;
      end
      8'b01100101 : begin
        _zz_wdata_3 = fifoDataBuffer_101;
      end
      8'b01100110 : begin
        _zz_wdata_3 = fifoDataBuffer_102;
      end
      8'b01100111 : begin
        _zz_wdata_3 = fifoDataBuffer_103;
      end
      8'b01101000 : begin
        _zz_wdata_3 = fifoDataBuffer_104;
      end
      8'b01101001 : begin
        _zz_wdata_3 = fifoDataBuffer_105;
      end
      8'b01101010 : begin
        _zz_wdata_3 = fifoDataBuffer_106;
      end
      8'b01101011 : begin
        _zz_wdata_3 = fifoDataBuffer_107;
      end
      8'b01101100 : begin
        _zz_wdata_3 = fifoDataBuffer_108;
      end
      8'b01101101 : begin
        _zz_wdata_3 = fifoDataBuffer_109;
      end
      8'b01101110 : begin
        _zz_wdata_3 = fifoDataBuffer_110;
      end
      8'b01101111 : begin
        _zz_wdata_3 = fifoDataBuffer_111;
      end
      8'b01110000 : begin
        _zz_wdata_3 = fifoDataBuffer_112;
      end
      8'b01110001 : begin
        _zz_wdata_3 = fifoDataBuffer_113;
      end
      8'b01110010 : begin
        _zz_wdata_3 = fifoDataBuffer_114;
      end
      8'b01110011 : begin
        _zz_wdata_3 = fifoDataBuffer_115;
      end
      8'b01110100 : begin
        _zz_wdata_3 = fifoDataBuffer_116;
      end
      8'b01110101 : begin
        _zz_wdata_3 = fifoDataBuffer_117;
      end
      8'b01110110 : begin
        _zz_wdata_3 = fifoDataBuffer_118;
      end
      8'b01110111 : begin
        _zz_wdata_3 = fifoDataBuffer_119;
      end
      8'b01111000 : begin
        _zz_wdata_3 = fifoDataBuffer_120;
      end
      8'b01111001 : begin
        _zz_wdata_3 = fifoDataBuffer_121;
      end
      8'b01111010 : begin
        _zz_wdata_3 = fifoDataBuffer_122;
      end
      8'b01111011 : begin
        _zz_wdata_3 = fifoDataBuffer_123;
      end
      8'b01111100 : begin
        _zz_wdata_3 = fifoDataBuffer_124;
      end
      8'b01111101 : begin
        _zz_wdata_3 = fifoDataBuffer_125;
      end
      8'b01111110 : begin
        _zz_wdata_3 = fifoDataBuffer_126;
      end
      8'b01111111 : begin
        _zz_wdata_3 = fifoDataBuffer_127;
      end
      8'b10000000 : begin
        _zz_wdata_3 = fifoDataBuffer_128;
      end
      8'b10000001 : begin
        _zz_wdata_3 = fifoDataBuffer_129;
      end
      8'b10000010 : begin
        _zz_wdata_3 = fifoDataBuffer_130;
      end
      8'b10000011 : begin
        _zz_wdata_3 = fifoDataBuffer_131;
      end
      8'b10000100 : begin
        _zz_wdata_3 = fifoDataBuffer_132;
      end
      8'b10000101 : begin
        _zz_wdata_3 = fifoDataBuffer_133;
      end
      8'b10000110 : begin
        _zz_wdata_3 = fifoDataBuffer_134;
      end
      8'b10000111 : begin
        _zz_wdata_3 = fifoDataBuffer_135;
      end
      8'b10001000 : begin
        _zz_wdata_3 = fifoDataBuffer_136;
      end
      8'b10001001 : begin
        _zz_wdata_3 = fifoDataBuffer_137;
      end
      8'b10001010 : begin
        _zz_wdata_3 = fifoDataBuffer_138;
      end
      8'b10001011 : begin
        _zz_wdata_3 = fifoDataBuffer_139;
      end
      8'b10001100 : begin
        _zz_wdata_3 = fifoDataBuffer_140;
      end
      8'b10001101 : begin
        _zz_wdata_3 = fifoDataBuffer_141;
      end
      8'b10001110 : begin
        _zz_wdata_3 = fifoDataBuffer_142;
      end
      8'b10001111 : begin
        _zz_wdata_3 = fifoDataBuffer_143;
      end
      8'b10010000 : begin
        _zz_wdata_3 = fifoDataBuffer_144;
      end
      8'b10010001 : begin
        _zz_wdata_3 = fifoDataBuffer_145;
      end
      8'b10010010 : begin
        _zz_wdata_3 = fifoDataBuffer_146;
      end
      8'b10010011 : begin
        _zz_wdata_3 = fifoDataBuffer_147;
      end
      8'b10010100 : begin
        _zz_wdata_3 = fifoDataBuffer_148;
      end
      8'b10010101 : begin
        _zz_wdata_3 = fifoDataBuffer_149;
      end
      8'b10010110 : begin
        _zz_wdata_3 = fifoDataBuffer_150;
      end
      8'b10010111 : begin
        _zz_wdata_3 = fifoDataBuffer_151;
      end
      8'b10011000 : begin
        _zz_wdata_3 = fifoDataBuffer_152;
      end
      8'b10011001 : begin
        _zz_wdata_3 = fifoDataBuffer_153;
      end
      8'b10011010 : begin
        _zz_wdata_3 = fifoDataBuffer_154;
      end
      8'b10011011 : begin
        _zz_wdata_3 = fifoDataBuffer_155;
      end
      8'b10011100 : begin
        _zz_wdata_3 = fifoDataBuffer_156;
      end
      8'b10011101 : begin
        _zz_wdata_3 = fifoDataBuffer_157;
      end
      8'b10011110 : begin
        _zz_wdata_3 = fifoDataBuffer_158;
      end
      8'b10011111 : begin
        _zz_wdata_3 = fifoDataBuffer_159;
      end
      8'b10100000 : begin
        _zz_wdata_3 = fifoDataBuffer_160;
      end
      8'b10100001 : begin
        _zz_wdata_3 = fifoDataBuffer_161;
      end
      8'b10100010 : begin
        _zz_wdata_3 = fifoDataBuffer_162;
      end
      8'b10100011 : begin
        _zz_wdata_3 = fifoDataBuffer_163;
      end
      8'b10100100 : begin
        _zz_wdata_3 = fifoDataBuffer_164;
      end
      8'b10100101 : begin
        _zz_wdata_3 = fifoDataBuffer_165;
      end
      8'b10100110 : begin
        _zz_wdata_3 = fifoDataBuffer_166;
      end
      8'b10100111 : begin
        _zz_wdata_3 = fifoDataBuffer_167;
      end
      8'b10101000 : begin
        _zz_wdata_3 = fifoDataBuffer_168;
      end
      8'b10101001 : begin
        _zz_wdata_3 = fifoDataBuffer_169;
      end
      8'b10101010 : begin
        _zz_wdata_3 = fifoDataBuffer_170;
      end
      8'b10101011 : begin
        _zz_wdata_3 = fifoDataBuffer_171;
      end
      8'b10101100 : begin
        _zz_wdata_3 = fifoDataBuffer_172;
      end
      8'b10101101 : begin
        _zz_wdata_3 = fifoDataBuffer_173;
      end
      8'b10101110 : begin
        _zz_wdata_3 = fifoDataBuffer_174;
      end
      8'b10101111 : begin
        _zz_wdata_3 = fifoDataBuffer_175;
      end
      8'b10110000 : begin
        _zz_wdata_3 = fifoDataBuffer_176;
      end
      8'b10110001 : begin
        _zz_wdata_3 = fifoDataBuffer_177;
      end
      8'b10110010 : begin
        _zz_wdata_3 = fifoDataBuffer_178;
      end
      8'b10110011 : begin
        _zz_wdata_3 = fifoDataBuffer_179;
      end
      8'b10110100 : begin
        _zz_wdata_3 = fifoDataBuffer_180;
      end
      8'b10110101 : begin
        _zz_wdata_3 = fifoDataBuffer_181;
      end
      8'b10110110 : begin
        _zz_wdata_3 = fifoDataBuffer_182;
      end
      8'b10110111 : begin
        _zz_wdata_3 = fifoDataBuffer_183;
      end
      8'b10111000 : begin
        _zz_wdata_3 = fifoDataBuffer_184;
      end
      8'b10111001 : begin
        _zz_wdata_3 = fifoDataBuffer_185;
      end
      8'b10111010 : begin
        _zz_wdata_3 = fifoDataBuffer_186;
      end
      8'b10111011 : begin
        _zz_wdata_3 = fifoDataBuffer_187;
      end
      8'b10111100 : begin
        _zz_wdata_3 = fifoDataBuffer_188;
      end
      8'b10111101 : begin
        _zz_wdata_3 = fifoDataBuffer_189;
      end
      8'b10111110 : begin
        _zz_wdata_3 = fifoDataBuffer_190;
      end
      8'b10111111 : begin
        _zz_wdata_3 = fifoDataBuffer_191;
      end
      8'b11000000 : begin
        _zz_wdata_3 = fifoDataBuffer_192;
      end
      8'b11000001 : begin
        _zz_wdata_3 = fifoDataBuffer_193;
      end
      8'b11000010 : begin
        _zz_wdata_3 = fifoDataBuffer_194;
      end
      8'b11000011 : begin
        _zz_wdata_3 = fifoDataBuffer_195;
      end
      8'b11000100 : begin
        _zz_wdata_3 = fifoDataBuffer_196;
      end
      8'b11000101 : begin
        _zz_wdata_3 = fifoDataBuffer_197;
      end
      8'b11000110 : begin
        _zz_wdata_3 = fifoDataBuffer_198;
      end
      8'b11000111 : begin
        _zz_wdata_3 = fifoDataBuffer_199;
      end
      8'b11001000 : begin
        _zz_wdata_3 = fifoDataBuffer_200;
      end
      8'b11001001 : begin
        _zz_wdata_3 = fifoDataBuffer_201;
      end
      8'b11001010 : begin
        _zz_wdata_3 = fifoDataBuffer_202;
      end
      8'b11001011 : begin
        _zz_wdata_3 = fifoDataBuffer_203;
      end
      8'b11001100 : begin
        _zz_wdata_3 = fifoDataBuffer_204;
      end
      8'b11001101 : begin
        _zz_wdata_3 = fifoDataBuffer_205;
      end
      8'b11001110 : begin
        _zz_wdata_3 = fifoDataBuffer_206;
      end
      8'b11001111 : begin
        _zz_wdata_3 = fifoDataBuffer_207;
      end
      8'b11010000 : begin
        _zz_wdata_3 = fifoDataBuffer_208;
      end
      8'b11010001 : begin
        _zz_wdata_3 = fifoDataBuffer_209;
      end
      8'b11010010 : begin
        _zz_wdata_3 = fifoDataBuffer_210;
      end
      8'b11010011 : begin
        _zz_wdata_3 = fifoDataBuffer_211;
      end
      8'b11010100 : begin
        _zz_wdata_3 = fifoDataBuffer_212;
      end
      8'b11010101 : begin
        _zz_wdata_3 = fifoDataBuffer_213;
      end
      8'b11010110 : begin
        _zz_wdata_3 = fifoDataBuffer_214;
      end
      8'b11010111 : begin
        _zz_wdata_3 = fifoDataBuffer_215;
      end
      8'b11011000 : begin
        _zz_wdata_3 = fifoDataBuffer_216;
      end
      8'b11011001 : begin
        _zz_wdata_3 = fifoDataBuffer_217;
      end
      8'b11011010 : begin
        _zz_wdata_3 = fifoDataBuffer_218;
      end
      8'b11011011 : begin
        _zz_wdata_3 = fifoDataBuffer_219;
      end
      8'b11011100 : begin
        _zz_wdata_3 = fifoDataBuffer_220;
      end
      8'b11011101 : begin
        _zz_wdata_3 = fifoDataBuffer_221;
      end
      8'b11011110 : begin
        _zz_wdata_3 = fifoDataBuffer_222;
      end
      8'b11011111 : begin
        _zz_wdata_3 = fifoDataBuffer_223;
      end
      8'b11100000 : begin
        _zz_wdata_3 = fifoDataBuffer_224;
      end
      8'b11100001 : begin
        _zz_wdata_3 = fifoDataBuffer_225;
      end
      8'b11100010 : begin
        _zz_wdata_3 = fifoDataBuffer_226;
      end
      8'b11100011 : begin
        _zz_wdata_3 = fifoDataBuffer_227;
      end
      8'b11100100 : begin
        _zz_wdata_3 = fifoDataBuffer_228;
      end
      8'b11100101 : begin
        _zz_wdata_3 = fifoDataBuffer_229;
      end
      8'b11100110 : begin
        _zz_wdata_3 = fifoDataBuffer_230;
      end
      8'b11100111 : begin
        _zz_wdata_3 = fifoDataBuffer_231;
      end
      8'b11101000 : begin
        _zz_wdata_3 = fifoDataBuffer_232;
      end
      8'b11101001 : begin
        _zz_wdata_3 = fifoDataBuffer_233;
      end
      8'b11101010 : begin
        _zz_wdata_3 = fifoDataBuffer_234;
      end
      8'b11101011 : begin
        _zz_wdata_3 = fifoDataBuffer_235;
      end
      8'b11101100 : begin
        _zz_wdata_3 = fifoDataBuffer_236;
      end
      8'b11101101 : begin
        _zz_wdata_3 = fifoDataBuffer_237;
      end
      8'b11101110 : begin
        _zz_wdata_3 = fifoDataBuffer_238;
      end
      8'b11101111 : begin
        _zz_wdata_3 = fifoDataBuffer_239;
      end
      8'b11110000 : begin
        _zz_wdata_3 = fifoDataBuffer_240;
      end
      8'b11110001 : begin
        _zz_wdata_3 = fifoDataBuffer_241;
      end
      8'b11110010 : begin
        _zz_wdata_3 = fifoDataBuffer_242;
      end
      8'b11110011 : begin
        _zz_wdata_3 = fifoDataBuffer_243;
      end
      8'b11110100 : begin
        _zz_wdata_3 = fifoDataBuffer_244;
      end
      8'b11110101 : begin
        _zz_wdata_3 = fifoDataBuffer_245;
      end
      8'b11110110 : begin
        _zz_wdata_3 = fifoDataBuffer_246;
      end
      8'b11110111 : begin
        _zz_wdata_3 = fifoDataBuffer_247;
      end
      8'b11111000 : begin
        _zz_wdata_3 = fifoDataBuffer_248;
      end
      8'b11111001 : begin
        _zz_wdata_3 = fifoDataBuffer_249;
      end
      8'b11111010 : begin
        _zz_wdata_3 = fifoDataBuffer_250;
      end
      8'b11111011 : begin
        _zz_wdata_3 = fifoDataBuffer_251;
      end
      8'b11111100 : begin
        _zz_wdata_3 = fifoDataBuffer_252;
      end
      8'b11111101 : begin
        _zz_wdata_3 = fifoDataBuffer_253;
      end
      8'b11111110 : begin
        _zz_wdata_3 = fifoDataBuffer_254;
      end
      default : begin
        _zz_wdata_3 = fifoDataBuffer_255;
      end
    endcase
  end

  always @(*) begin
    _zz_wdata = 1'b0;
    if(when_Axi4WriteMaster_l118) begin
      _zz_wdata = 1'b1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(_zz_when_Axi4WriteMaster_l61) begin
      _zz_1 = 1'b1;
    end
  end

  assign _zz_when_Axi4WriteMaster_l61 = (_zz_wdata_2 == 9'h100);
  assign _zz_2 = (_zz_when_Axi4WriteMaster_l61 && _zz_wdata);
  always @(*) begin
    if(_zz_2) begin
      _zz_wdata_1 = 9'h0;
    end else begin
      _zz_wdata_1 = (_zz_wdata_2 + _zz__zz_wdata_1);
    end
    if(_zz_1) begin
      _zz_wdata_1 = 9'h0;
    end
  end

  always @(*) begin
    _zz_when_Axi4WriteMaster_l53 = 1'b0;
    if(when_Axi4WriteMaster_l47) begin
      _zz_when_Axi4WriteMaster_l53 = 1'b1;
    end
  end

  always @(*) begin
    _zz_3 = 1'b0;
    if(when_Axi4WriteMaster_l61) begin
      _zz_3 = 1'b1;
    end
  end

  assign _zz_when_Axi4WriteMaster_l53_3 = (_zz_when_Axi4WriteMaster_l53_2 == 9'h100);
  assign _zz_4 = (_zz_when_Axi4WriteMaster_l53_3 && _zz_when_Axi4WriteMaster_l53);
  always @(*) begin
    if(_zz_4) begin
      _zz_when_Axi4WriteMaster_l53_1 = 9'h0;
    end else begin
      _zz_when_Axi4WriteMaster_l53_1 = (_zz_when_Axi4WriteMaster_l53_2 + _zz__zz_when_Axi4WriteMaster_l53_1);
    end
    if(_zz_3) begin
      _zz_when_Axi4WriteMaster_l53_1 = 9'h0;
    end
  end

  assign when_Axi4WriteMaster_l47 = (fifoValid && fifoReady);
  assign _zz_5 = ({255'd0,1'b1} <<< _zz__zz_5);
  always @(*) begin
    fifoReady = 1'b0;
    if(when_Axi4WriteMaster_l53) begin
      fifoReady = 1'b1;
    end
  end

  assign when_Axi4WriteMaster_l53 = (! _zz_when_Axi4WriteMaster_l53_3);
  assign when_Axi4WriteMaster_l61 = (_zz_when_Axi4WriteMaster_l61 && (bresp == 2'b00));
  assign when_Axi4WriteMaster_l70 = (awValid && awReady);
  assign Axi4Incr_validSize = awsize[1 : 0];
  assign Axi4Incr_highCat = axi4Interface_address[31 : 12];
  assign Axi4Incr_sizeValue = {(2'b10 == Axi4Incr_validSize),{(2'b01 == Axi4Incr_validSize),(2'b00 == Axi4Incr_validSize)}};
  assign Axi4Incr_alignMask = {10'd0, _zz_Axi4Incr_alignMask};
  assign Axi4Incr_base = (_zz_Axi4Incr_base & (~ Axi4Incr_alignMask));
  assign Axi4Incr_baseIncr = (Axi4Incr_base + _zz_Axi4Incr_baseIncr);
  always @(*) begin
    casez(awlen)
      8'b????1??? : begin
        _zz_Axi4Incr_wrapCase = 2'b11;
      end
      8'b?????1?? : begin
        _zz_Axi4Incr_wrapCase = 2'b10;
      end
      8'b??????1? : begin
        _zz_Axi4Incr_wrapCase = 2'b01;
      end
      default : begin
        _zz_Axi4Incr_wrapCase = 2'b00;
      end
    endcase
  end

  assign Axi4Incr_wrapCase = (_zz_Axi4Incr_wrapCase_1 + _zz_Axi4Incr_wrapCase_2);
  always @(*) begin
    case(awburst)
      2'b00 : begin
        Axi4Incr_result = axi4Interface_address;
      end
      2'b10 : begin
        Axi4Incr_result = {Axi4Incr_highCat,_zz_Axi4Incr_result};
      end
      default : begin
        Axi4Incr_result = {Axi4Incr_highCat,Axi4Incr_baseIncr};
      end
    endcase
  end

  assign awValid = wValid;
  assign when_Axi4WriteMaster_l87 = (_zz_wdata_2 == 9'h0);
  always @(*) begin
    if(_zz_when_Axi4WriteMaster_l61) begin
      awaddr = axi4Interface_address;
    end else begin
      awaddr = axi4Interface_initialAddress;
    end
  end

  assign awid = 1'b0;
  assign awregion = 4'b0000;
  assign awburst = 2'b01;
  assign awlen = 8'hff;
  assign awsize = 3'b100;
  assign awlock = 1'b0;
  assign awcache = 4'b0000;
  assign awqos = 4'b0000;
  assign awprot = 3'b000;
  always @(*) begin
    wdata = 32'h0;
    if(wValid) begin
      wdata = _zz_wdata_3;
    end
  end

  assign when_Axi4WriteMaster_l118 = (wValid && wReady);
  always @(*) begin
    wValid = 1'b0;
    if(when_Axi4WriteMaster_l124) begin
      wValid = 1'b1;
    end
  end

  assign when_Axi4WriteMaster_l124 = ((9'h0 < _zz_when_Axi4WriteMaster_l53_2) && (! _zz_when_Axi4WriteMaster_l61));
  assign wstrb = 4'b1111;
  assign wlast = (_zz_wdata_2 == 9'h0ff);
  assign bReady = 1'b0;
  assign araddr = 32'h0;
  assign arid = 1'b0;
  assign arregion = 4'b0000;
  assign arburst = 2'b01;
  assign arlen = 8'hff;
  assign arsize = 3'b100;
  assign arlock = 1'b0;
  assign arcache = 4'b0000;
  assign arqos = 4'b0000;
  assign arprot = 3'b000;
  assign arValid = 1'b0;
  assign rReady = 1'b0;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _zz_wdata_2 <= 9'h0;
      _zz_when_Axi4WriteMaster_l53_2 <= 9'h0;
      fifoDataBuffer_0 <= 32'h0;
      fifoDataBuffer_1 <= 32'h0;
      fifoDataBuffer_2 <= 32'h0;
      fifoDataBuffer_3 <= 32'h0;
      fifoDataBuffer_4 <= 32'h0;
      fifoDataBuffer_5 <= 32'h0;
      fifoDataBuffer_6 <= 32'h0;
      fifoDataBuffer_7 <= 32'h0;
      fifoDataBuffer_8 <= 32'h0;
      fifoDataBuffer_9 <= 32'h0;
      fifoDataBuffer_10 <= 32'h0;
      fifoDataBuffer_11 <= 32'h0;
      fifoDataBuffer_12 <= 32'h0;
      fifoDataBuffer_13 <= 32'h0;
      fifoDataBuffer_14 <= 32'h0;
      fifoDataBuffer_15 <= 32'h0;
      fifoDataBuffer_16 <= 32'h0;
      fifoDataBuffer_17 <= 32'h0;
      fifoDataBuffer_18 <= 32'h0;
      fifoDataBuffer_19 <= 32'h0;
      fifoDataBuffer_20 <= 32'h0;
      fifoDataBuffer_21 <= 32'h0;
      fifoDataBuffer_22 <= 32'h0;
      fifoDataBuffer_23 <= 32'h0;
      fifoDataBuffer_24 <= 32'h0;
      fifoDataBuffer_25 <= 32'h0;
      fifoDataBuffer_26 <= 32'h0;
      fifoDataBuffer_27 <= 32'h0;
      fifoDataBuffer_28 <= 32'h0;
      fifoDataBuffer_29 <= 32'h0;
      fifoDataBuffer_30 <= 32'h0;
      fifoDataBuffer_31 <= 32'h0;
      fifoDataBuffer_32 <= 32'h0;
      fifoDataBuffer_33 <= 32'h0;
      fifoDataBuffer_34 <= 32'h0;
      fifoDataBuffer_35 <= 32'h0;
      fifoDataBuffer_36 <= 32'h0;
      fifoDataBuffer_37 <= 32'h0;
      fifoDataBuffer_38 <= 32'h0;
      fifoDataBuffer_39 <= 32'h0;
      fifoDataBuffer_40 <= 32'h0;
      fifoDataBuffer_41 <= 32'h0;
      fifoDataBuffer_42 <= 32'h0;
      fifoDataBuffer_43 <= 32'h0;
      fifoDataBuffer_44 <= 32'h0;
      fifoDataBuffer_45 <= 32'h0;
      fifoDataBuffer_46 <= 32'h0;
      fifoDataBuffer_47 <= 32'h0;
      fifoDataBuffer_48 <= 32'h0;
      fifoDataBuffer_49 <= 32'h0;
      fifoDataBuffer_50 <= 32'h0;
      fifoDataBuffer_51 <= 32'h0;
      fifoDataBuffer_52 <= 32'h0;
      fifoDataBuffer_53 <= 32'h0;
      fifoDataBuffer_54 <= 32'h0;
      fifoDataBuffer_55 <= 32'h0;
      fifoDataBuffer_56 <= 32'h0;
      fifoDataBuffer_57 <= 32'h0;
      fifoDataBuffer_58 <= 32'h0;
      fifoDataBuffer_59 <= 32'h0;
      fifoDataBuffer_60 <= 32'h0;
      fifoDataBuffer_61 <= 32'h0;
      fifoDataBuffer_62 <= 32'h0;
      fifoDataBuffer_63 <= 32'h0;
      fifoDataBuffer_64 <= 32'h0;
      fifoDataBuffer_65 <= 32'h0;
      fifoDataBuffer_66 <= 32'h0;
      fifoDataBuffer_67 <= 32'h0;
      fifoDataBuffer_68 <= 32'h0;
      fifoDataBuffer_69 <= 32'h0;
      fifoDataBuffer_70 <= 32'h0;
      fifoDataBuffer_71 <= 32'h0;
      fifoDataBuffer_72 <= 32'h0;
      fifoDataBuffer_73 <= 32'h0;
      fifoDataBuffer_74 <= 32'h0;
      fifoDataBuffer_75 <= 32'h0;
      fifoDataBuffer_76 <= 32'h0;
      fifoDataBuffer_77 <= 32'h0;
      fifoDataBuffer_78 <= 32'h0;
      fifoDataBuffer_79 <= 32'h0;
      fifoDataBuffer_80 <= 32'h0;
      fifoDataBuffer_81 <= 32'h0;
      fifoDataBuffer_82 <= 32'h0;
      fifoDataBuffer_83 <= 32'h0;
      fifoDataBuffer_84 <= 32'h0;
      fifoDataBuffer_85 <= 32'h0;
      fifoDataBuffer_86 <= 32'h0;
      fifoDataBuffer_87 <= 32'h0;
      fifoDataBuffer_88 <= 32'h0;
      fifoDataBuffer_89 <= 32'h0;
      fifoDataBuffer_90 <= 32'h0;
      fifoDataBuffer_91 <= 32'h0;
      fifoDataBuffer_92 <= 32'h0;
      fifoDataBuffer_93 <= 32'h0;
      fifoDataBuffer_94 <= 32'h0;
      fifoDataBuffer_95 <= 32'h0;
      fifoDataBuffer_96 <= 32'h0;
      fifoDataBuffer_97 <= 32'h0;
      fifoDataBuffer_98 <= 32'h0;
      fifoDataBuffer_99 <= 32'h0;
      fifoDataBuffer_100 <= 32'h0;
      fifoDataBuffer_101 <= 32'h0;
      fifoDataBuffer_102 <= 32'h0;
      fifoDataBuffer_103 <= 32'h0;
      fifoDataBuffer_104 <= 32'h0;
      fifoDataBuffer_105 <= 32'h0;
      fifoDataBuffer_106 <= 32'h0;
      fifoDataBuffer_107 <= 32'h0;
      fifoDataBuffer_108 <= 32'h0;
      fifoDataBuffer_109 <= 32'h0;
      fifoDataBuffer_110 <= 32'h0;
      fifoDataBuffer_111 <= 32'h0;
      fifoDataBuffer_112 <= 32'h0;
      fifoDataBuffer_113 <= 32'h0;
      fifoDataBuffer_114 <= 32'h0;
      fifoDataBuffer_115 <= 32'h0;
      fifoDataBuffer_116 <= 32'h0;
      fifoDataBuffer_117 <= 32'h0;
      fifoDataBuffer_118 <= 32'h0;
      fifoDataBuffer_119 <= 32'h0;
      fifoDataBuffer_120 <= 32'h0;
      fifoDataBuffer_121 <= 32'h0;
      fifoDataBuffer_122 <= 32'h0;
      fifoDataBuffer_123 <= 32'h0;
      fifoDataBuffer_124 <= 32'h0;
      fifoDataBuffer_125 <= 32'h0;
      fifoDataBuffer_126 <= 32'h0;
      fifoDataBuffer_127 <= 32'h0;
      fifoDataBuffer_128 <= 32'h0;
      fifoDataBuffer_129 <= 32'h0;
      fifoDataBuffer_130 <= 32'h0;
      fifoDataBuffer_131 <= 32'h0;
      fifoDataBuffer_132 <= 32'h0;
      fifoDataBuffer_133 <= 32'h0;
      fifoDataBuffer_134 <= 32'h0;
      fifoDataBuffer_135 <= 32'h0;
      fifoDataBuffer_136 <= 32'h0;
      fifoDataBuffer_137 <= 32'h0;
      fifoDataBuffer_138 <= 32'h0;
      fifoDataBuffer_139 <= 32'h0;
      fifoDataBuffer_140 <= 32'h0;
      fifoDataBuffer_141 <= 32'h0;
      fifoDataBuffer_142 <= 32'h0;
      fifoDataBuffer_143 <= 32'h0;
      fifoDataBuffer_144 <= 32'h0;
      fifoDataBuffer_145 <= 32'h0;
      fifoDataBuffer_146 <= 32'h0;
      fifoDataBuffer_147 <= 32'h0;
      fifoDataBuffer_148 <= 32'h0;
      fifoDataBuffer_149 <= 32'h0;
      fifoDataBuffer_150 <= 32'h0;
      fifoDataBuffer_151 <= 32'h0;
      fifoDataBuffer_152 <= 32'h0;
      fifoDataBuffer_153 <= 32'h0;
      fifoDataBuffer_154 <= 32'h0;
      fifoDataBuffer_155 <= 32'h0;
      fifoDataBuffer_156 <= 32'h0;
      fifoDataBuffer_157 <= 32'h0;
      fifoDataBuffer_158 <= 32'h0;
      fifoDataBuffer_159 <= 32'h0;
      fifoDataBuffer_160 <= 32'h0;
      fifoDataBuffer_161 <= 32'h0;
      fifoDataBuffer_162 <= 32'h0;
      fifoDataBuffer_163 <= 32'h0;
      fifoDataBuffer_164 <= 32'h0;
      fifoDataBuffer_165 <= 32'h0;
      fifoDataBuffer_166 <= 32'h0;
      fifoDataBuffer_167 <= 32'h0;
      fifoDataBuffer_168 <= 32'h0;
      fifoDataBuffer_169 <= 32'h0;
      fifoDataBuffer_170 <= 32'h0;
      fifoDataBuffer_171 <= 32'h0;
      fifoDataBuffer_172 <= 32'h0;
      fifoDataBuffer_173 <= 32'h0;
      fifoDataBuffer_174 <= 32'h0;
      fifoDataBuffer_175 <= 32'h0;
      fifoDataBuffer_176 <= 32'h0;
      fifoDataBuffer_177 <= 32'h0;
      fifoDataBuffer_178 <= 32'h0;
      fifoDataBuffer_179 <= 32'h0;
      fifoDataBuffer_180 <= 32'h0;
      fifoDataBuffer_181 <= 32'h0;
      fifoDataBuffer_182 <= 32'h0;
      fifoDataBuffer_183 <= 32'h0;
      fifoDataBuffer_184 <= 32'h0;
      fifoDataBuffer_185 <= 32'h0;
      fifoDataBuffer_186 <= 32'h0;
      fifoDataBuffer_187 <= 32'h0;
      fifoDataBuffer_188 <= 32'h0;
      fifoDataBuffer_189 <= 32'h0;
      fifoDataBuffer_190 <= 32'h0;
      fifoDataBuffer_191 <= 32'h0;
      fifoDataBuffer_192 <= 32'h0;
      fifoDataBuffer_193 <= 32'h0;
      fifoDataBuffer_194 <= 32'h0;
      fifoDataBuffer_195 <= 32'h0;
      fifoDataBuffer_196 <= 32'h0;
      fifoDataBuffer_197 <= 32'h0;
      fifoDataBuffer_198 <= 32'h0;
      fifoDataBuffer_199 <= 32'h0;
      fifoDataBuffer_200 <= 32'h0;
      fifoDataBuffer_201 <= 32'h0;
      fifoDataBuffer_202 <= 32'h0;
      fifoDataBuffer_203 <= 32'h0;
      fifoDataBuffer_204 <= 32'h0;
      fifoDataBuffer_205 <= 32'h0;
      fifoDataBuffer_206 <= 32'h0;
      fifoDataBuffer_207 <= 32'h0;
      fifoDataBuffer_208 <= 32'h0;
      fifoDataBuffer_209 <= 32'h0;
      fifoDataBuffer_210 <= 32'h0;
      fifoDataBuffer_211 <= 32'h0;
      fifoDataBuffer_212 <= 32'h0;
      fifoDataBuffer_213 <= 32'h0;
      fifoDataBuffer_214 <= 32'h0;
      fifoDataBuffer_215 <= 32'h0;
      fifoDataBuffer_216 <= 32'h0;
      fifoDataBuffer_217 <= 32'h0;
      fifoDataBuffer_218 <= 32'h0;
      fifoDataBuffer_219 <= 32'h0;
      fifoDataBuffer_220 <= 32'h0;
      fifoDataBuffer_221 <= 32'h0;
      fifoDataBuffer_222 <= 32'h0;
      fifoDataBuffer_223 <= 32'h0;
      fifoDataBuffer_224 <= 32'h0;
      fifoDataBuffer_225 <= 32'h0;
      fifoDataBuffer_226 <= 32'h0;
      fifoDataBuffer_227 <= 32'h0;
      fifoDataBuffer_228 <= 32'h0;
      fifoDataBuffer_229 <= 32'h0;
      fifoDataBuffer_230 <= 32'h0;
      fifoDataBuffer_231 <= 32'h0;
      fifoDataBuffer_232 <= 32'h0;
      fifoDataBuffer_233 <= 32'h0;
      fifoDataBuffer_234 <= 32'h0;
      fifoDataBuffer_235 <= 32'h0;
      fifoDataBuffer_236 <= 32'h0;
      fifoDataBuffer_237 <= 32'h0;
      fifoDataBuffer_238 <= 32'h0;
      fifoDataBuffer_239 <= 32'h0;
      fifoDataBuffer_240 <= 32'h0;
      fifoDataBuffer_241 <= 32'h0;
      fifoDataBuffer_242 <= 32'h0;
      fifoDataBuffer_243 <= 32'h0;
      fifoDataBuffer_244 <= 32'h0;
      fifoDataBuffer_245 <= 32'h0;
      fifoDataBuffer_246 <= 32'h0;
      fifoDataBuffer_247 <= 32'h0;
      fifoDataBuffer_248 <= 32'h0;
      fifoDataBuffer_249 <= 32'h0;
      fifoDataBuffer_250 <= 32'h0;
      fifoDataBuffer_251 <= 32'h0;
      fifoDataBuffer_252 <= 32'h0;
      fifoDataBuffer_253 <= 32'h0;
      fifoDataBuffer_254 <= 32'h0;
      fifoDataBuffer_255 <= 32'h0;
      axi4Interface_address <= 32'h0;
      axi4Interface_initialAddress <= 32'h0;
    end else begin
      _zz_wdata_2 <= _zz_wdata_1;
      _zz_when_Axi4WriteMaster_l53_2 <= _zz_when_Axi4WriteMaster_l53_1;
      if(when_Axi4WriteMaster_l47) begin
        if(_zz_5[0]) begin
          fifoDataBuffer_0 <= fifoPayload;
        end
        if(_zz_5[1]) begin
          fifoDataBuffer_1 <= fifoPayload;
        end
        if(_zz_5[2]) begin
          fifoDataBuffer_2 <= fifoPayload;
        end
        if(_zz_5[3]) begin
          fifoDataBuffer_3 <= fifoPayload;
        end
        if(_zz_5[4]) begin
          fifoDataBuffer_4 <= fifoPayload;
        end
        if(_zz_5[5]) begin
          fifoDataBuffer_5 <= fifoPayload;
        end
        if(_zz_5[6]) begin
          fifoDataBuffer_6 <= fifoPayload;
        end
        if(_zz_5[7]) begin
          fifoDataBuffer_7 <= fifoPayload;
        end
        if(_zz_5[8]) begin
          fifoDataBuffer_8 <= fifoPayload;
        end
        if(_zz_5[9]) begin
          fifoDataBuffer_9 <= fifoPayload;
        end
        if(_zz_5[10]) begin
          fifoDataBuffer_10 <= fifoPayload;
        end
        if(_zz_5[11]) begin
          fifoDataBuffer_11 <= fifoPayload;
        end
        if(_zz_5[12]) begin
          fifoDataBuffer_12 <= fifoPayload;
        end
        if(_zz_5[13]) begin
          fifoDataBuffer_13 <= fifoPayload;
        end
        if(_zz_5[14]) begin
          fifoDataBuffer_14 <= fifoPayload;
        end
        if(_zz_5[15]) begin
          fifoDataBuffer_15 <= fifoPayload;
        end
        if(_zz_5[16]) begin
          fifoDataBuffer_16 <= fifoPayload;
        end
        if(_zz_5[17]) begin
          fifoDataBuffer_17 <= fifoPayload;
        end
        if(_zz_5[18]) begin
          fifoDataBuffer_18 <= fifoPayload;
        end
        if(_zz_5[19]) begin
          fifoDataBuffer_19 <= fifoPayload;
        end
        if(_zz_5[20]) begin
          fifoDataBuffer_20 <= fifoPayload;
        end
        if(_zz_5[21]) begin
          fifoDataBuffer_21 <= fifoPayload;
        end
        if(_zz_5[22]) begin
          fifoDataBuffer_22 <= fifoPayload;
        end
        if(_zz_5[23]) begin
          fifoDataBuffer_23 <= fifoPayload;
        end
        if(_zz_5[24]) begin
          fifoDataBuffer_24 <= fifoPayload;
        end
        if(_zz_5[25]) begin
          fifoDataBuffer_25 <= fifoPayload;
        end
        if(_zz_5[26]) begin
          fifoDataBuffer_26 <= fifoPayload;
        end
        if(_zz_5[27]) begin
          fifoDataBuffer_27 <= fifoPayload;
        end
        if(_zz_5[28]) begin
          fifoDataBuffer_28 <= fifoPayload;
        end
        if(_zz_5[29]) begin
          fifoDataBuffer_29 <= fifoPayload;
        end
        if(_zz_5[30]) begin
          fifoDataBuffer_30 <= fifoPayload;
        end
        if(_zz_5[31]) begin
          fifoDataBuffer_31 <= fifoPayload;
        end
        if(_zz_5[32]) begin
          fifoDataBuffer_32 <= fifoPayload;
        end
        if(_zz_5[33]) begin
          fifoDataBuffer_33 <= fifoPayload;
        end
        if(_zz_5[34]) begin
          fifoDataBuffer_34 <= fifoPayload;
        end
        if(_zz_5[35]) begin
          fifoDataBuffer_35 <= fifoPayload;
        end
        if(_zz_5[36]) begin
          fifoDataBuffer_36 <= fifoPayload;
        end
        if(_zz_5[37]) begin
          fifoDataBuffer_37 <= fifoPayload;
        end
        if(_zz_5[38]) begin
          fifoDataBuffer_38 <= fifoPayload;
        end
        if(_zz_5[39]) begin
          fifoDataBuffer_39 <= fifoPayload;
        end
        if(_zz_5[40]) begin
          fifoDataBuffer_40 <= fifoPayload;
        end
        if(_zz_5[41]) begin
          fifoDataBuffer_41 <= fifoPayload;
        end
        if(_zz_5[42]) begin
          fifoDataBuffer_42 <= fifoPayload;
        end
        if(_zz_5[43]) begin
          fifoDataBuffer_43 <= fifoPayload;
        end
        if(_zz_5[44]) begin
          fifoDataBuffer_44 <= fifoPayload;
        end
        if(_zz_5[45]) begin
          fifoDataBuffer_45 <= fifoPayload;
        end
        if(_zz_5[46]) begin
          fifoDataBuffer_46 <= fifoPayload;
        end
        if(_zz_5[47]) begin
          fifoDataBuffer_47 <= fifoPayload;
        end
        if(_zz_5[48]) begin
          fifoDataBuffer_48 <= fifoPayload;
        end
        if(_zz_5[49]) begin
          fifoDataBuffer_49 <= fifoPayload;
        end
        if(_zz_5[50]) begin
          fifoDataBuffer_50 <= fifoPayload;
        end
        if(_zz_5[51]) begin
          fifoDataBuffer_51 <= fifoPayload;
        end
        if(_zz_5[52]) begin
          fifoDataBuffer_52 <= fifoPayload;
        end
        if(_zz_5[53]) begin
          fifoDataBuffer_53 <= fifoPayload;
        end
        if(_zz_5[54]) begin
          fifoDataBuffer_54 <= fifoPayload;
        end
        if(_zz_5[55]) begin
          fifoDataBuffer_55 <= fifoPayload;
        end
        if(_zz_5[56]) begin
          fifoDataBuffer_56 <= fifoPayload;
        end
        if(_zz_5[57]) begin
          fifoDataBuffer_57 <= fifoPayload;
        end
        if(_zz_5[58]) begin
          fifoDataBuffer_58 <= fifoPayload;
        end
        if(_zz_5[59]) begin
          fifoDataBuffer_59 <= fifoPayload;
        end
        if(_zz_5[60]) begin
          fifoDataBuffer_60 <= fifoPayload;
        end
        if(_zz_5[61]) begin
          fifoDataBuffer_61 <= fifoPayload;
        end
        if(_zz_5[62]) begin
          fifoDataBuffer_62 <= fifoPayload;
        end
        if(_zz_5[63]) begin
          fifoDataBuffer_63 <= fifoPayload;
        end
        if(_zz_5[64]) begin
          fifoDataBuffer_64 <= fifoPayload;
        end
        if(_zz_5[65]) begin
          fifoDataBuffer_65 <= fifoPayload;
        end
        if(_zz_5[66]) begin
          fifoDataBuffer_66 <= fifoPayload;
        end
        if(_zz_5[67]) begin
          fifoDataBuffer_67 <= fifoPayload;
        end
        if(_zz_5[68]) begin
          fifoDataBuffer_68 <= fifoPayload;
        end
        if(_zz_5[69]) begin
          fifoDataBuffer_69 <= fifoPayload;
        end
        if(_zz_5[70]) begin
          fifoDataBuffer_70 <= fifoPayload;
        end
        if(_zz_5[71]) begin
          fifoDataBuffer_71 <= fifoPayload;
        end
        if(_zz_5[72]) begin
          fifoDataBuffer_72 <= fifoPayload;
        end
        if(_zz_5[73]) begin
          fifoDataBuffer_73 <= fifoPayload;
        end
        if(_zz_5[74]) begin
          fifoDataBuffer_74 <= fifoPayload;
        end
        if(_zz_5[75]) begin
          fifoDataBuffer_75 <= fifoPayload;
        end
        if(_zz_5[76]) begin
          fifoDataBuffer_76 <= fifoPayload;
        end
        if(_zz_5[77]) begin
          fifoDataBuffer_77 <= fifoPayload;
        end
        if(_zz_5[78]) begin
          fifoDataBuffer_78 <= fifoPayload;
        end
        if(_zz_5[79]) begin
          fifoDataBuffer_79 <= fifoPayload;
        end
        if(_zz_5[80]) begin
          fifoDataBuffer_80 <= fifoPayload;
        end
        if(_zz_5[81]) begin
          fifoDataBuffer_81 <= fifoPayload;
        end
        if(_zz_5[82]) begin
          fifoDataBuffer_82 <= fifoPayload;
        end
        if(_zz_5[83]) begin
          fifoDataBuffer_83 <= fifoPayload;
        end
        if(_zz_5[84]) begin
          fifoDataBuffer_84 <= fifoPayload;
        end
        if(_zz_5[85]) begin
          fifoDataBuffer_85 <= fifoPayload;
        end
        if(_zz_5[86]) begin
          fifoDataBuffer_86 <= fifoPayload;
        end
        if(_zz_5[87]) begin
          fifoDataBuffer_87 <= fifoPayload;
        end
        if(_zz_5[88]) begin
          fifoDataBuffer_88 <= fifoPayload;
        end
        if(_zz_5[89]) begin
          fifoDataBuffer_89 <= fifoPayload;
        end
        if(_zz_5[90]) begin
          fifoDataBuffer_90 <= fifoPayload;
        end
        if(_zz_5[91]) begin
          fifoDataBuffer_91 <= fifoPayload;
        end
        if(_zz_5[92]) begin
          fifoDataBuffer_92 <= fifoPayload;
        end
        if(_zz_5[93]) begin
          fifoDataBuffer_93 <= fifoPayload;
        end
        if(_zz_5[94]) begin
          fifoDataBuffer_94 <= fifoPayload;
        end
        if(_zz_5[95]) begin
          fifoDataBuffer_95 <= fifoPayload;
        end
        if(_zz_5[96]) begin
          fifoDataBuffer_96 <= fifoPayload;
        end
        if(_zz_5[97]) begin
          fifoDataBuffer_97 <= fifoPayload;
        end
        if(_zz_5[98]) begin
          fifoDataBuffer_98 <= fifoPayload;
        end
        if(_zz_5[99]) begin
          fifoDataBuffer_99 <= fifoPayload;
        end
        if(_zz_5[100]) begin
          fifoDataBuffer_100 <= fifoPayload;
        end
        if(_zz_5[101]) begin
          fifoDataBuffer_101 <= fifoPayload;
        end
        if(_zz_5[102]) begin
          fifoDataBuffer_102 <= fifoPayload;
        end
        if(_zz_5[103]) begin
          fifoDataBuffer_103 <= fifoPayload;
        end
        if(_zz_5[104]) begin
          fifoDataBuffer_104 <= fifoPayload;
        end
        if(_zz_5[105]) begin
          fifoDataBuffer_105 <= fifoPayload;
        end
        if(_zz_5[106]) begin
          fifoDataBuffer_106 <= fifoPayload;
        end
        if(_zz_5[107]) begin
          fifoDataBuffer_107 <= fifoPayload;
        end
        if(_zz_5[108]) begin
          fifoDataBuffer_108 <= fifoPayload;
        end
        if(_zz_5[109]) begin
          fifoDataBuffer_109 <= fifoPayload;
        end
        if(_zz_5[110]) begin
          fifoDataBuffer_110 <= fifoPayload;
        end
        if(_zz_5[111]) begin
          fifoDataBuffer_111 <= fifoPayload;
        end
        if(_zz_5[112]) begin
          fifoDataBuffer_112 <= fifoPayload;
        end
        if(_zz_5[113]) begin
          fifoDataBuffer_113 <= fifoPayload;
        end
        if(_zz_5[114]) begin
          fifoDataBuffer_114 <= fifoPayload;
        end
        if(_zz_5[115]) begin
          fifoDataBuffer_115 <= fifoPayload;
        end
        if(_zz_5[116]) begin
          fifoDataBuffer_116 <= fifoPayload;
        end
        if(_zz_5[117]) begin
          fifoDataBuffer_117 <= fifoPayload;
        end
        if(_zz_5[118]) begin
          fifoDataBuffer_118 <= fifoPayload;
        end
        if(_zz_5[119]) begin
          fifoDataBuffer_119 <= fifoPayload;
        end
        if(_zz_5[120]) begin
          fifoDataBuffer_120 <= fifoPayload;
        end
        if(_zz_5[121]) begin
          fifoDataBuffer_121 <= fifoPayload;
        end
        if(_zz_5[122]) begin
          fifoDataBuffer_122 <= fifoPayload;
        end
        if(_zz_5[123]) begin
          fifoDataBuffer_123 <= fifoPayload;
        end
        if(_zz_5[124]) begin
          fifoDataBuffer_124 <= fifoPayload;
        end
        if(_zz_5[125]) begin
          fifoDataBuffer_125 <= fifoPayload;
        end
        if(_zz_5[126]) begin
          fifoDataBuffer_126 <= fifoPayload;
        end
        if(_zz_5[127]) begin
          fifoDataBuffer_127 <= fifoPayload;
        end
        if(_zz_5[128]) begin
          fifoDataBuffer_128 <= fifoPayload;
        end
        if(_zz_5[129]) begin
          fifoDataBuffer_129 <= fifoPayload;
        end
        if(_zz_5[130]) begin
          fifoDataBuffer_130 <= fifoPayload;
        end
        if(_zz_5[131]) begin
          fifoDataBuffer_131 <= fifoPayload;
        end
        if(_zz_5[132]) begin
          fifoDataBuffer_132 <= fifoPayload;
        end
        if(_zz_5[133]) begin
          fifoDataBuffer_133 <= fifoPayload;
        end
        if(_zz_5[134]) begin
          fifoDataBuffer_134 <= fifoPayload;
        end
        if(_zz_5[135]) begin
          fifoDataBuffer_135 <= fifoPayload;
        end
        if(_zz_5[136]) begin
          fifoDataBuffer_136 <= fifoPayload;
        end
        if(_zz_5[137]) begin
          fifoDataBuffer_137 <= fifoPayload;
        end
        if(_zz_5[138]) begin
          fifoDataBuffer_138 <= fifoPayload;
        end
        if(_zz_5[139]) begin
          fifoDataBuffer_139 <= fifoPayload;
        end
        if(_zz_5[140]) begin
          fifoDataBuffer_140 <= fifoPayload;
        end
        if(_zz_5[141]) begin
          fifoDataBuffer_141 <= fifoPayload;
        end
        if(_zz_5[142]) begin
          fifoDataBuffer_142 <= fifoPayload;
        end
        if(_zz_5[143]) begin
          fifoDataBuffer_143 <= fifoPayload;
        end
        if(_zz_5[144]) begin
          fifoDataBuffer_144 <= fifoPayload;
        end
        if(_zz_5[145]) begin
          fifoDataBuffer_145 <= fifoPayload;
        end
        if(_zz_5[146]) begin
          fifoDataBuffer_146 <= fifoPayload;
        end
        if(_zz_5[147]) begin
          fifoDataBuffer_147 <= fifoPayload;
        end
        if(_zz_5[148]) begin
          fifoDataBuffer_148 <= fifoPayload;
        end
        if(_zz_5[149]) begin
          fifoDataBuffer_149 <= fifoPayload;
        end
        if(_zz_5[150]) begin
          fifoDataBuffer_150 <= fifoPayload;
        end
        if(_zz_5[151]) begin
          fifoDataBuffer_151 <= fifoPayload;
        end
        if(_zz_5[152]) begin
          fifoDataBuffer_152 <= fifoPayload;
        end
        if(_zz_5[153]) begin
          fifoDataBuffer_153 <= fifoPayload;
        end
        if(_zz_5[154]) begin
          fifoDataBuffer_154 <= fifoPayload;
        end
        if(_zz_5[155]) begin
          fifoDataBuffer_155 <= fifoPayload;
        end
        if(_zz_5[156]) begin
          fifoDataBuffer_156 <= fifoPayload;
        end
        if(_zz_5[157]) begin
          fifoDataBuffer_157 <= fifoPayload;
        end
        if(_zz_5[158]) begin
          fifoDataBuffer_158 <= fifoPayload;
        end
        if(_zz_5[159]) begin
          fifoDataBuffer_159 <= fifoPayload;
        end
        if(_zz_5[160]) begin
          fifoDataBuffer_160 <= fifoPayload;
        end
        if(_zz_5[161]) begin
          fifoDataBuffer_161 <= fifoPayload;
        end
        if(_zz_5[162]) begin
          fifoDataBuffer_162 <= fifoPayload;
        end
        if(_zz_5[163]) begin
          fifoDataBuffer_163 <= fifoPayload;
        end
        if(_zz_5[164]) begin
          fifoDataBuffer_164 <= fifoPayload;
        end
        if(_zz_5[165]) begin
          fifoDataBuffer_165 <= fifoPayload;
        end
        if(_zz_5[166]) begin
          fifoDataBuffer_166 <= fifoPayload;
        end
        if(_zz_5[167]) begin
          fifoDataBuffer_167 <= fifoPayload;
        end
        if(_zz_5[168]) begin
          fifoDataBuffer_168 <= fifoPayload;
        end
        if(_zz_5[169]) begin
          fifoDataBuffer_169 <= fifoPayload;
        end
        if(_zz_5[170]) begin
          fifoDataBuffer_170 <= fifoPayload;
        end
        if(_zz_5[171]) begin
          fifoDataBuffer_171 <= fifoPayload;
        end
        if(_zz_5[172]) begin
          fifoDataBuffer_172 <= fifoPayload;
        end
        if(_zz_5[173]) begin
          fifoDataBuffer_173 <= fifoPayload;
        end
        if(_zz_5[174]) begin
          fifoDataBuffer_174 <= fifoPayload;
        end
        if(_zz_5[175]) begin
          fifoDataBuffer_175 <= fifoPayload;
        end
        if(_zz_5[176]) begin
          fifoDataBuffer_176 <= fifoPayload;
        end
        if(_zz_5[177]) begin
          fifoDataBuffer_177 <= fifoPayload;
        end
        if(_zz_5[178]) begin
          fifoDataBuffer_178 <= fifoPayload;
        end
        if(_zz_5[179]) begin
          fifoDataBuffer_179 <= fifoPayload;
        end
        if(_zz_5[180]) begin
          fifoDataBuffer_180 <= fifoPayload;
        end
        if(_zz_5[181]) begin
          fifoDataBuffer_181 <= fifoPayload;
        end
        if(_zz_5[182]) begin
          fifoDataBuffer_182 <= fifoPayload;
        end
        if(_zz_5[183]) begin
          fifoDataBuffer_183 <= fifoPayload;
        end
        if(_zz_5[184]) begin
          fifoDataBuffer_184 <= fifoPayload;
        end
        if(_zz_5[185]) begin
          fifoDataBuffer_185 <= fifoPayload;
        end
        if(_zz_5[186]) begin
          fifoDataBuffer_186 <= fifoPayload;
        end
        if(_zz_5[187]) begin
          fifoDataBuffer_187 <= fifoPayload;
        end
        if(_zz_5[188]) begin
          fifoDataBuffer_188 <= fifoPayload;
        end
        if(_zz_5[189]) begin
          fifoDataBuffer_189 <= fifoPayload;
        end
        if(_zz_5[190]) begin
          fifoDataBuffer_190 <= fifoPayload;
        end
        if(_zz_5[191]) begin
          fifoDataBuffer_191 <= fifoPayload;
        end
        if(_zz_5[192]) begin
          fifoDataBuffer_192 <= fifoPayload;
        end
        if(_zz_5[193]) begin
          fifoDataBuffer_193 <= fifoPayload;
        end
        if(_zz_5[194]) begin
          fifoDataBuffer_194 <= fifoPayload;
        end
        if(_zz_5[195]) begin
          fifoDataBuffer_195 <= fifoPayload;
        end
        if(_zz_5[196]) begin
          fifoDataBuffer_196 <= fifoPayload;
        end
        if(_zz_5[197]) begin
          fifoDataBuffer_197 <= fifoPayload;
        end
        if(_zz_5[198]) begin
          fifoDataBuffer_198 <= fifoPayload;
        end
        if(_zz_5[199]) begin
          fifoDataBuffer_199 <= fifoPayload;
        end
        if(_zz_5[200]) begin
          fifoDataBuffer_200 <= fifoPayload;
        end
        if(_zz_5[201]) begin
          fifoDataBuffer_201 <= fifoPayload;
        end
        if(_zz_5[202]) begin
          fifoDataBuffer_202 <= fifoPayload;
        end
        if(_zz_5[203]) begin
          fifoDataBuffer_203 <= fifoPayload;
        end
        if(_zz_5[204]) begin
          fifoDataBuffer_204 <= fifoPayload;
        end
        if(_zz_5[205]) begin
          fifoDataBuffer_205 <= fifoPayload;
        end
        if(_zz_5[206]) begin
          fifoDataBuffer_206 <= fifoPayload;
        end
        if(_zz_5[207]) begin
          fifoDataBuffer_207 <= fifoPayload;
        end
        if(_zz_5[208]) begin
          fifoDataBuffer_208 <= fifoPayload;
        end
        if(_zz_5[209]) begin
          fifoDataBuffer_209 <= fifoPayload;
        end
        if(_zz_5[210]) begin
          fifoDataBuffer_210 <= fifoPayload;
        end
        if(_zz_5[211]) begin
          fifoDataBuffer_211 <= fifoPayload;
        end
        if(_zz_5[212]) begin
          fifoDataBuffer_212 <= fifoPayload;
        end
        if(_zz_5[213]) begin
          fifoDataBuffer_213 <= fifoPayload;
        end
        if(_zz_5[214]) begin
          fifoDataBuffer_214 <= fifoPayload;
        end
        if(_zz_5[215]) begin
          fifoDataBuffer_215 <= fifoPayload;
        end
        if(_zz_5[216]) begin
          fifoDataBuffer_216 <= fifoPayload;
        end
        if(_zz_5[217]) begin
          fifoDataBuffer_217 <= fifoPayload;
        end
        if(_zz_5[218]) begin
          fifoDataBuffer_218 <= fifoPayload;
        end
        if(_zz_5[219]) begin
          fifoDataBuffer_219 <= fifoPayload;
        end
        if(_zz_5[220]) begin
          fifoDataBuffer_220 <= fifoPayload;
        end
        if(_zz_5[221]) begin
          fifoDataBuffer_221 <= fifoPayload;
        end
        if(_zz_5[222]) begin
          fifoDataBuffer_222 <= fifoPayload;
        end
        if(_zz_5[223]) begin
          fifoDataBuffer_223 <= fifoPayload;
        end
        if(_zz_5[224]) begin
          fifoDataBuffer_224 <= fifoPayload;
        end
        if(_zz_5[225]) begin
          fifoDataBuffer_225 <= fifoPayload;
        end
        if(_zz_5[226]) begin
          fifoDataBuffer_226 <= fifoPayload;
        end
        if(_zz_5[227]) begin
          fifoDataBuffer_227 <= fifoPayload;
        end
        if(_zz_5[228]) begin
          fifoDataBuffer_228 <= fifoPayload;
        end
        if(_zz_5[229]) begin
          fifoDataBuffer_229 <= fifoPayload;
        end
        if(_zz_5[230]) begin
          fifoDataBuffer_230 <= fifoPayload;
        end
        if(_zz_5[231]) begin
          fifoDataBuffer_231 <= fifoPayload;
        end
        if(_zz_5[232]) begin
          fifoDataBuffer_232 <= fifoPayload;
        end
        if(_zz_5[233]) begin
          fifoDataBuffer_233 <= fifoPayload;
        end
        if(_zz_5[234]) begin
          fifoDataBuffer_234 <= fifoPayload;
        end
        if(_zz_5[235]) begin
          fifoDataBuffer_235 <= fifoPayload;
        end
        if(_zz_5[236]) begin
          fifoDataBuffer_236 <= fifoPayload;
        end
        if(_zz_5[237]) begin
          fifoDataBuffer_237 <= fifoPayload;
        end
        if(_zz_5[238]) begin
          fifoDataBuffer_238 <= fifoPayload;
        end
        if(_zz_5[239]) begin
          fifoDataBuffer_239 <= fifoPayload;
        end
        if(_zz_5[240]) begin
          fifoDataBuffer_240 <= fifoPayload;
        end
        if(_zz_5[241]) begin
          fifoDataBuffer_241 <= fifoPayload;
        end
        if(_zz_5[242]) begin
          fifoDataBuffer_242 <= fifoPayload;
        end
        if(_zz_5[243]) begin
          fifoDataBuffer_243 <= fifoPayload;
        end
        if(_zz_5[244]) begin
          fifoDataBuffer_244 <= fifoPayload;
        end
        if(_zz_5[245]) begin
          fifoDataBuffer_245 <= fifoPayload;
        end
        if(_zz_5[246]) begin
          fifoDataBuffer_246 <= fifoPayload;
        end
        if(_zz_5[247]) begin
          fifoDataBuffer_247 <= fifoPayload;
        end
        if(_zz_5[248]) begin
          fifoDataBuffer_248 <= fifoPayload;
        end
        if(_zz_5[249]) begin
          fifoDataBuffer_249 <= fifoPayload;
        end
        if(_zz_5[250]) begin
          fifoDataBuffer_250 <= fifoPayload;
        end
        if(_zz_5[251]) begin
          fifoDataBuffer_251 <= fifoPayload;
        end
        if(_zz_5[252]) begin
          fifoDataBuffer_252 <= fifoPayload;
        end
        if(_zz_5[253]) begin
          fifoDataBuffer_253 <= fifoPayload;
        end
        if(_zz_5[254]) begin
          fifoDataBuffer_254 <= fifoPayload;
        end
        if(_zz_5[255]) begin
          fifoDataBuffer_255 <= fifoPayload;
        end
      end
      if(when_Axi4WriteMaster_l70) begin
        axi4Interface_address <= Axi4Incr_result;
      end
      if(when_Axi4WriteMaster_l87) begin
        axi4Interface_initialAddress <= axi4Interface_address;
      end
    end
  end


endmodule
