// Generator : SpinalHDL v1.6.1    git head : 3bf789d53b1b5a36974196e2d591342e15ddf28c
// Component : arraySlice
// Git hash  : c0a2a0d076879a33f43d275808257504bfb7d141

`timescale 1ns/1ps 

module arraySlice (
  input               inputStreamArrayData_valid,
  output reg          inputStreamArrayData_ready,
  input      [31:0]   inputStreamArrayData_payload,
  input      [5:0]    inputFeatureMapWidth,
  input      [5:0]    inputFeatureMapHeight,
  input      [2:0]    outputFeatureMapHeight,
  input      [2:0]    outputFeatureMapWidth,
  output reg          outputStreamArrayData_0_valid,
  input               outputStreamArrayData_0_ready,
  output reg [31:0]   outputStreamArrayData_0_payload,
  output reg          outputStreamArrayData_1_valid,
  input               outputStreamArrayData_1_ready,
  output reg [31:0]   outputStreamArrayData_1_payload,
  output reg          outputStreamArrayData_2_valid,
  input               outputStreamArrayData_2_ready,
  output reg [31:0]   outputStreamArrayData_2_payload,
  output reg          outputStreamArrayData_3_valid,
  input               outputStreamArrayData_3_ready,
  output reg [31:0]   outputStreamArrayData_3_payload,
  output reg          outputStreamArrayData_4_valid,
  input               outputStreamArrayData_4_ready,
  output reg [31:0]   outputStreamArrayData_4_payload,
  output reg          outputStreamArrayData_5_valid,
  input               outputStreamArrayData_5_ready,
  output reg [31:0]   outputStreamArrayData_5_payload,
  output reg          outputStreamArrayData_6_valid,
  input               outputStreamArrayData_6_ready,
  output reg [31:0]   outputStreamArrayData_6_payload,
  output reg          outputStreamArrayData_7_valid,
  input               outputStreamArrayData_7_ready,
  output reg [31:0]   outputStreamArrayData_7_payload,
  input               clk,
  input               resetn
);
  localparam arraySliceStateMachine_enumDef_BOOT = 2'd0;
  localparam arraySliceStateMachine_enumDef_writeDataOnly = 2'd1;
  localparam arraySliceStateMachine_enumDef_readDataOnly = 2'd2;
  localparam arraySliceStateMachine_enumDef_readWriteData = 2'd3;

  reg                 fifoGroup_0_io_push_valid;
  reg        [31:0]   fifoGroup_0_io_push_payload;
  reg                 fifoGroup_0_io_pop_ready;
  reg                 fifoGroup_1_io_push_valid;
  reg        [31:0]   fifoGroup_1_io_push_payload;
  reg                 fifoGroup_1_io_pop_ready;
  reg                 fifoGroup_2_io_push_valid;
  reg        [31:0]   fifoGroup_2_io_push_payload;
  reg                 fifoGroup_2_io_pop_ready;
  reg                 fifoGroup_3_io_push_valid;
  reg        [31:0]   fifoGroup_3_io_push_payload;
  reg                 fifoGroup_3_io_pop_ready;
  reg                 fifoGroup_4_io_push_valid;
  reg        [31:0]   fifoGroup_4_io_push_payload;
  reg                 fifoGroup_4_io_pop_ready;
  reg                 fifoGroup_5_io_push_valid;
  reg        [31:0]   fifoGroup_5_io_push_payload;
  reg                 fifoGroup_5_io_pop_ready;
  reg                 fifoGroup_6_io_push_valid;
  reg        [31:0]   fifoGroup_6_io_push_payload;
  reg                 fifoGroup_6_io_pop_ready;
  reg                 fifoGroup_7_io_push_valid;
  reg        [31:0]   fifoGroup_7_io_push_payload;
  reg                 fifoGroup_7_io_pop_ready;
  reg                 fifoGroup_8_io_push_valid;
  reg        [31:0]   fifoGroup_8_io_push_payload;
  reg                 fifoGroup_8_io_pop_ready;
  reg                 fifoGroup_9_io_push_valid;
  reg        [31:0]   fifoGroup_9_io_push_payload;
  reg                 fifoGroup_9_io_pop_ready;
  reg                 fifoGroup_10_io_push_valid;
  reg        [31:0]   fifoGroup_10_io_push_payload;
  reg                 fifoGroup_10_io_pop_ready;
  reg                 fifoGroup_11_io_push_valid;
  reg        [31:0]   fifoGroup_11_io_push_payload;
  reg                 fifoGroup_11_io_pop_ready;
  reg                 fifoGroup_12_io_push_valid;
  reg        [31:0]   fifoGroup_12_io_push_payload;
  reg                 fifoGroup_12_io_pop_ready;
  reg                 fifoGroup_13_io_push_valid;
  reg        [31:0]   fifoGroup_13_io_push_payload;
  reg                 fifoGroup_13_io_pop_ready;
  reg                 fifoGroup_14_io_push_valid;
  reg        [31:0]   fifoGroup_14_io_push_payload;
  reg                 fifoGroup_14_io_pop_ready;
  reg                 fifoGroup_15_io_push_valid;
  reg        [31:0]   fifoGroup_15_io_push_payload;
  reg                 fifoGroup_15_io_pop_ready;
  reg                 fifoGroup_16_io_push_valid;
  reg        [31:0]   fifoGroup_16_io_push_payload;
  reg                 fifoGroup_16_io_pop_ready;
  reg                 fifoGroup_17_io_push_valid;
  reg        [31:0]   fifoGroup_17_io_push_payload;
  reg                 fifoGroup_17_io_pop_ready;
  reg                 fifoGroup_18_io_push_valid;
  reg        [31:0]   fifoGroup_18_io_push_payload;
  reg                 fifoGroup_18_io_pop_ready;
  reg                 fifoGroup_19_io_push_valid;
  reg        [31:0]   fifoGroup_19_io_push_payload;
  reg                 fifoGroup_19_io_pop_ready;
  reg                 fifoGroup_20_io_push_valid;
  reg        [31:0]   fifoGroup_20_io_push_payload;
  reg                 fifoGroup_20_io_pop_ready;
  reg                 fifoGroup_21_io_push_valid;
  reg        [31:0]   fifoGroup_21_io_push_payload;
  reg                 fifoGroup_21_io_pop_ready;
  reg                 fifoGroup_22_io_push_valid;
  reg        [31:0]   fifoGroup_22_io_push_payload;
  reg                 fifoGroup_22_io_pop_ready;
  reg                 fifoGroup_23_io_push_valid;
  reg        [31:0]   fifoGroup_23_io_push_payload;
  reg                 fifoGroup_23_io_pop_ready;
  reg                 fifoGroup_24_io_push_valid;
  reg        [31:0]   fifoGroup_24_io_push_payload;
  reg                 fifoGroup_24_io_pop_ready;
  reg                 fifoGroup_25_io_push_valid;
  reg        [31:0]   fifoGroup_25_io_push_payload;
  reg                 fifoGroup_25_io_pop_ready;
  reg                 fifoGroup_26_io_push_valid;
  reg        [31:0]   fifoGroup_26_io_push_payload;
  reg                 fifoGroup_26_io_pop_ready;
  reg                 fifoGroup_27_io_push_valid;
  reg        [31:0]   fifoGroup_27_io_push_payload;
  reg                 fifoGroup_27_io_pop_ready;
  reg                 fifoGroup_28_io_push_valid;
  reg        [31:0]   fifoGroup_28_io_push_payload;
  reg                 fifoGroup_28_io_pop_ready;
  reg                 fifoGroup_29_io_push_valid;
  reg        [31:0]   fifoGroup_29_io_push_payload;
  reg                 fifoGroup_29_io_pop_ready;
  reg                 fifoGroup_30_io_push_valid;
  reg        [31:0]   fifoGroup_30_io_push_payload;
  reg                 fifoGroup_30_io_pop_ready;
  reg                 fifoGroup_31_io_push_valid;
  reg        [31:0]   fifoGroup_31_io_push_payload;
  reg                 fifoGroup_31_io_pop_ready;
  reg                 fifoGroup_32_io_push_valid;
  reg        [31:0]   fifoGroup_32_io_push_payload;
  reg                 fifoGroup_32_io_pop_ready;
  reg                 fifoGroup_33_io_push_valid;
  reg        [31:0]   fifoGroup_33_io_push_payload;
  reg                 fifoGroup_33_io_pop_ready;
  reg                 fifoGroup_34_io_push_valid;
  reg        [31:0]   fifoGroup_34_io_push_payload;
  reg                 fifoGroup_34_io_pop_ready;
  reg                 fifoGroup_35_io_push_valid;
  reg        [31:0]   fifoGroup_35_io_push_payload;
  reg                 fifoGroup_35_io_pop_ready;
  reg                 fifoGroup_36_io_push_valid;
  reg        [31:0]   fifoGroup_36_io_push_payload;
  reg                 fifoGroup_36_io_pop_ready;
  reg                 fifoGroup_37_io_push_valid;
  reg        [31:0]   fifoGroup_37_io_push_payload;
  reg                 fifoGroup_37_io_pop_ready;
  reg                 fifoGroup_38_io_push_valid;
  reg        [31:0]   fifoGroup_38_io_push_payload;
  reg                 fifoGroup_38_io_pop_ready;
  reg                 fifoGroup_39_io_push_valid;
  reg        [31:0]   fifoGroup_39_io_push_payload;
  reg                 fifoGroup_39_io_pop_ready;
  reg                 fifoGroup_40_io_push_valid;
  reg        [31:0]   fifoGroup_40_io_push_payload;
  reg                 fifoGroup_40_io_pop_ready;
  reg                 fifoGroup_41_io_push_valid;
  reg        [31:0]   fifoGroup_41_io_push_payload;
  reg                 fifoGroup_41_io_pop_ready;
  reg                 fifoGroup_42_io_push_valid;
  reg        [31:0]   fifoGroup_42_io_push_payload;
  reg                 fifoGroup_42_io_pop_ready;
  reg                 fifoGroup_43_io_push_valid;
  reg        [31:0]   fifoGroup_43_io_push_payload;
  reg                 fifoGroup_43_io_pop_ready;
  reg                 fifoGroup_44_io_push_valid;
  reg        [31:0]   fifoGroup_44_io_push_payload;
  reg                 fifoGroup_44_io_pop_ready;
  reg                 fifoGroup_45_io_push_valid;
  reg        [31:0]   fifoGroup_45_io_push_payload;
  reg                 fifoGroup_45_io_pop_ready;
  reg                 fifoGroup_46_io_push_valid;
  reg        [31:0]   fifoGroup_46_io_push_payload;
  reg                 fifoGroup_46_io_pop_ready;
  reg                 fifoGroup_47_io_push_valid;
  reg        [31:0]   fifoGroup_47_io_push_payload;
  reg                 fifoGroup_47_io_pop_ready;
  reg                 fifoGroup_48_io_push_valid;
  reg        [31:0]   fifoGroup_48_io_push_payload;
  reg                 fifoGroup_48_io_pop_ready;
  reg                 fifoGroup_49_io_push_valid;
  reg        [31:0]   fifoGroup_49_io_push_payload;
  reg                 fifoGroup_49_io_pop_ready;
  reg                 fifoGroup_50_io_push_valid;
  reg        [31:0]   fifoGroup_50_io_push_payload;
  reg                 fifoGroup_50_io_pop_ready;
  reg                 fifoGroup_51_io_push_valid;
  reg        [31:0]   fifoGroup_51_io_push_payload;
  reg                 fifoGroup_51_io_pop_ready;
  reg                 fifoGroup_52_io_push_valid;
  reg        [31:0]   fifoGroup_52_io_push_payload;
  reg                 fifoGroup_52_io_pop_ready;
  reg                 fifoGroup_53_io_push_valid;
  reg        [31:0]   fifoGroup_53_io_push_payload;
  reg                 fifoGroup_53_io_pop_ready;
  reg                 fifoGroup_54_io_push_valid;
  reg        [31:0]   fifoGroup_54_io_push_payload;
  reg                 fifoGroup_54_io_pop_ready;
  reg                 fifoGroup_55_io_push_valid;
  reg        [31:0]   fifoGroup_55_io_push_payload;
  reg                 fifoGroup_55_io_pop_ready;
  reg                 fifoGroup_56_io_push_valid;
  reg        [31:0]   fifoGroup_56_io_push_payload;
  reg                 fifoGroup_56_io_pop_ready;
  reg                 fifoGroup_57_io_push_valid;
  reg        [31:0]   fifoGroup_57_io_push_payload;
  reg                 fifoGroup_57_io_pop_ready;
  reg                 fifoGroup_58_io_push_valid;
  reg        [31:0]   fifoGroup_58_io_push_payload;
  reg                 fifoGroup_58_io_pop_ready;
  reg                 fifoGroup_59_io_push_valid;
  reg        [31:0]   fifoGroup_59_io_push_payload;
  reg                 fifoGroup_59_io_pop_ready;
  reg                 fifoGroup_60_io_push_valid;
  reg        [31:0]   fifoGroup_60_io_push_payload;
  reg                 fifoGroup_60_io_pop_ready;
  reg                 fifoGroup_61_io_push_valid;
  reg        [31:0]   fifoGroup_61_io_push_payload;
  reg                 fifoGroup_61_io_pop_ready;
  reg                 fifoGroup_62_io_push_valid;
  reg        [31:0]   fifoGroup_62_io_push_payload;
  reg                 fifoGroup_62_io_pop_ready;
  reg                 fifoGroup_63_io_push_valid;
  reg        [31:0]   fifoGroup_63_io_push_payload;
  reg                 fifoGroup_63_io_pop_ready;
  wire                fifoGroup_0_io_push_ready;
  wire                fifoGroup_0_io_pop_valid;
  wire       [31:0]   fifoGroup_0_io_pop_payload;
  wire       [6:0]    fifoGroup_0_io_occupancy;
  wire       [6:0]    fifoGroup_0_io_availability;
  wire                fifoGroup_1_io_push_ready;
  wire                fifoGroup_1_io_pop_valid;
  wire       [31:0]   fifoGroup_1_io_pop_payload;
  wire       [6:0]    fifoGroup_1_io_occupancy;
  wire       [6:0]    fifoGroup_1_io_availability;
  wire                fifoGroup_2_io_push_ready;
  wire                fifoGroup_2_io_pop_valid;
  wire       [31:0]   fifoGroup_2_io_pop_payload;
  wire       [6:0]    fifoGroup_2_io_occupancy;
  wire       [6:0]    fifoGroup_2_io_availability;
  wire                fifoGroup_3_io_push_ready;
  wire                fifoGroup_3_io_pop_valid;
  wire       [31:0]   fifoGroup_3_io_pop_payload;
  wire       [6:0]    fifoGroup_3_io_occupancy;
  wire       [6:0]    fifoGroup_3_io_availability;
  wire                fifoGroup_4_io_push_ready;
  wire                fifoGroup_4_io_pop_valid;
  wire       [31:0]   fifoGroup_4_io_pop_payload;
  wire       [6:0]    fifoGroup_4_io_occupancy;
  wire       [6:0]    fifoGroup_4_io_availability;
  wire                fifoGroup_5_io_push_ready;
  wire                fifoGroup_5_io_pop_valid;
  wire       [31:0]   fifoGroup_5_io_pop_payload;
  wire       [6:0]    fifoGroup_5_io_occupancy;
  wire       [6:0]    fifoGroup_5_io_availability;
  wire                fifoGroup_6_io_push_ready;
  wire                fifoGroup_6_io_pop_valid;
  wire       [31:0]   fifoGroup_6_io_pop_payload;
  wire       [6:0]    fifoGroup_6_io_occupancy;
  wire       [6:0]    fifoGroup_6_io_availability;
  wire                fifoGroup_7_io_push_ready;
  wire                fifoGroup_7_io_pop_valid;
  wire       [31:0]   fifoGroup_7_io_pop_payload;
  wire       [6:0]    fifoGroup_7_io_occupancy;
  wire       [6:0]    fifoGroup_7_io_availability;
  wire                fifoGroup_8_io_push_ready;
  wire                fifoGroup_8_io_pop_valid;
  wire       [31:0]   fifoGroup_8_io_pop_payload;
  wire       [6:0]    fifoGroup_8_io_occupancy;
  wire       [6:0]    fifoGroup_8_io_availability;
  wire                fifoGroup_9_io_push_ready;
  wire                fifoGroup_9_io_pop_valid;
  wire       [31:0]   fifoGroup_9_io_pop_payload;
  wire       [6:0]    fifoGroup_9_io_occupancy;
  wire       [6:0]    fifoGroup_9_io_availability;
  wire                fifoGroup_10_io_push_ready;
  wire                fifoGroup_10_io_pop_valid;
  wire       [31:0]   fifoGroup_10_io_pop_payload;
  wire       [6:0]    fifoGroup_10_io_occupancy;
  wire       [6:0]    fifoGroup_10_io_availability;
  wire                fifoGroup_11_io_push_ready;
  wire                fifoGroup_11_io_pop_valid;
  wire       [31:0]   fifoGroup_11_io_pop_payload;
  wire       [6:0]    fifoGroup_11_io_occupancy;
  wire       [6:0]    fifoGroup_11_io_availability;
  wire                fifoGroup_12_io_push_ready;
  wire                fifoGroup_12_io_pop_valid;
  wire       [31:0]   fifoGroup_12_io_pop_payload;
  wire       [6:0]    fifoGroup_12_io_occupancy;
  wire       [6:0]    fifoGroup_12_io_availability;
  wire                fifoGroup_13_io_push_ready;
  wire                fifoGroup_13_io_pop_valid;
  wire       [31:0]   fifoGroup_13_io_pop_payload;
  wire       [6:0]    fifoGroup_13_io_occupancy;
  wire       [6:0]    fifoGroup_13_io_availability;
  wire                fifoGroup_14_io_push_ready;
  wire                fifoGroup_14_io_pop_valid;
  wire       [31:0]   fifoGroup_14_io_pop_payload;
  wire       [6:0]    fifoGroup_14_io_occupancy;
  wire       [6:0]    fifoGroup_14_io_availability;
  wire                fifoGroup_15_io_push_ready;
  wire                fifoGroup_15_io_pop_valid;
  wire       [31:0]   fifoGroup_15_io_pop_payload;
  wire       [6:0]    fifoGroup_15_io_occupancy;
  wire       [6:0]    fifoGroup_15_io_availability;
  wire                fifoGroup_16_io_push_ready;
  wire                fifoGroup_16_io_pop_valid;
  wire       [31:0]   fifoGroup_16_io_pop_payload;
  wire       [6:0]    fifoGroup_16_io_occupancy;
  wire       [6:0]    fifoGroup_16_io_availability;
  wire                fifoGroup_17_io_push_ready;
  wire                fifoGroup_17_io_pop_valid;
  wire       [31:0]   fifoGroup_17_io_pop_payload;
  wire       [6:0]    fifoGroup_17_io_occupancy;
  wire       [6:0]    fifoGroup_17_io_availability;
  wire                fifoGroup_18_io_push_ready;
  wire                fifoGroup_18_io_pop_valid;
  wire       [31:0]   fifoGroup_18_io_pop_payload;
  wire       [6:0]    fifoGroup_18_io_occupancy;
  wire       [6:0]    fifoGroup_18_io_availability;
  wire                fifoGroup_19_io_push_ready;
  wire                fifoGroup_19_io_pop_valid;
  wire       [31:0]   fifoGroup_19_io_pop_payload;
  wire       [6:0]    fifoGroup_19_io_occupancy;
  wire       [6:0]    fifoGroup_19_io_availability;
  wire                fifoGroup_20_io_push_ready;
  wire                fifoGroup_20_io_pop_valid;
  wire       [31:0]   fifoGroup_20_io_pop_payload;
  wire       [6:0]    fifoGroup_20_io_occupancy;
  wire       [6:0]    fifoGroup_20_io_availability;
  wire                fifoGroup_21_io_push_ready;
  wire                fifoGroup_21_io_pop_valid;
  wire       [31:0]   fifoGroup_21_io_pop_payload;
  wire       [6:0]    fifoGroup_21_io_occupancy;
  wire       [6:0]    fifoGroup_21_io_availability;
  wire                fifoGroup_22_io_push_ready;
  wire                fifoGroup_22_io_pop_valid;
  wire       [31:0]   fifoGroup_22_io_pop_payload;
  wire       [6:0]    fifoGroup_22_io_occupancy;
  wire       [6:0]    fifoGroup_22_io_availability;
  wire                fifoGroup_23_io_push_ready;
  wire                fifoGroup_23_io_pop_valid;
  wire       [31:0]   fifoGroup_23_io_pop_payload;
  wire       [6:0]    fifoGroup_23_io_occupancy;
  wire       [6:0]    fifoGroup_23_io_availability;
  wire                fifoGroup_24_io_push_ready;
  wire                fifoGroup_24_io_pop_valid;
  wire       [31:0]   fifoGroup_24_io_pop_payload;
  wire       [6:0]    fifoGroup_24_io_occupancy;
  wire       [6:0]    fifoGroup_24_io_availability;
  wire                fifoGroup_25_io_push_ready;
  wire                fifoGroup_25_io_pop_valid;
  wire       [31:0]   fifoGroup_25_io_pop_payload;
  wire       [6:0]    fifoGroup_25_io_occupancy;
  wire       [6:0]    fifoGroup_25_io_availability;
  wire                fifoGroup_26_io_push_ready;
  wire                fifoGroup_26_io_pop_valid;
  wire       [31:0]   fifoGroup_26_io_pop_payload;
  wire       [6:0]    fifoGroup_26_io_occupancy;
  wire       [6:0]    fifoGroup_26_io_availability;
  wire                fifoGroup_27_io_push_ready;
  wire                fifoGroup_27_io_pop_valid;
  wire       [31:0]   fifoGroup_27_io_pop_payload;
  wire       [6:0]    fifoGroup_27_io_occupancy;
  wire       [6:0]    fifoGroup_27_io_availability;
  wire                fifoGroup_28_io_push_ready;
  wire                fifoGroup_28_io_pop_valid;
  wire       [31:0]   fifoGroup_28_io_pop_payload;
  wire       [6:0]    fifoGroup_28_io_occupancy;
  wire       [6:0]    fifoGroup_28_io_availability;
  wire                fifoGroup_29_io_push_ready;
  wire                fifoGroup_29_io_pop_valid;
  wire       [31:0]   fifoGroup_29_io_pop_payload;
  wire       [6:0]    fifoGroup_29_io_occupancy;
  wire       [6:0]    fifoGroup_29_io_availability;
  wire                fifoGroup_30_io_push_ready;
  wire                fifoGroup_30_io_pop_valid;
  wire       [31:0]   fifoGroup_30_io_pop_payload;
  wire       [6:0]    fifoGroup_30_io_occupancy;
  wire       [6:0]    fifoGroup_30_io_availability;
  wire                fifoGroup_31_io_push_ready;
  wire                fifoGroup_31_io_pop_valid;
  wire       [31:0]   fifoGroup_31_io_pop_payload;
  wire       [6:0]    fifoGroup_31_io_occupancy;
  wire       [6:0]    fifoGroup_31_io_availability;
  wire                fifoGroup_32_io_push_ready;
  wire                fifoGroup_32_io_pop_valid;
  wire       [31:0]   fifoGroup_32_io_pop_payload;
  wire       [6:0]    fifoGroup_32_io_occupancy;
  wire       [6:0]    fifoGroup_32_io_availability;
  wire                fifoGroup_33_io_push_ready;
  wire                fifoGroup_33_io_pop_valid;
  wire       [31:0]   fifoGroup_33_io_pop_payload;
  wire       [6:0]    fifoGroup_33_io_occupancy;
  wire       [6:0]    fifoGroup_33_io_availability;
  wire                fifoGroup_34_io_push_ready;
  wire                fifoGroup_34_io_pop_valid;
  wire       [31:0]   fifoGroup_34_io_pop_payload;
  wire       [6:0]    fifoGroup_34_io_occupancy;
  wire       [6:0]    fifoGroup_34_io_availability;
  wire                fifoGroup_35_io_push_ready;
  wire                fifoGroup_35_io_pop_valid;
  wire       [31:0]   fifoGroup_35_io_pop_payload;
  wire       [6:0]    fifoGroup_35_io_occupancy;
  wire       [6:0]    fifoGroup_35_io_availability;
  wire                fifoGroup_36_io_push_ready;
  wire                fifoGroup_36_io_pop_valid;
  wire       [31:0]   fifoGroup_36_io_pop_payload;
  wire       [6:0]    fifoGroup_36_io_occupancy;
  wire       [6:0]    fifoGroup_36_io_availability;
  wire                fifoGroup_37_io_push_ready;
  wire                fifoGroup_37_io_pop_valid;
  wire       [31:0]   fifoGroup_37_io_pop_payload;
  wire       [6:0]    fifoGroup_37_io_occupancy;
  wire       [6:0]    fifoGroup_37_io_availability;
  wire                fifoGroup_38_io_push_ready;
  wire                fifoGroup_38_io_pop_valid;
  wire       [31:0]   fifoGroup_38_io_pop_payload;
  wire       [6:0]    fifoGroup_38_io_occupancy;
  wire       [6:0]    fifoGroup_38_io_availability;
  wire                fifoGroup_39_io_push_ready;
  wire                fifoGroup_39_io_pop_valid;
  wire       [31:0]   fifoGroup_39_io_pop_payload;
  wire       [6:0]    fifoGroup_39_io_occupancy;
  wire       [6:0]    fifoGroup_39_io_availability;
  wire                fifoGroup_40_io_push_ready;
  wire                fifoGroup_40_io_pop_valid;
  wire       [31:0]   fifoGroup_40_io_pop_payload;
  wire       [6:0]    fifoGroup_40_io_occupancy;
  wire       [6:0]    fifoGroup_40_io_availability;
  wire                fifoGroup_41_io_push_ready;
  wire                fifoGroup_41_io_pop_valid;
  wire       [31:0]   fifoGroup_41_io_pop_payload;
  wire       [6:0]    fifoGroup_41_io_occupancy;
  wire       [6:0]    fifoGroup_41_io_availability;
  wire                fifoGroup_42_io_push_ready;
  wire                fifoGroup_42_io_pop_valid;
  wire       [31:0]   fifoGroup_42_io_pop_payload;
  wire       [6:0]    fifoGroup_42_io_occupancy;
  wire       [6:0]    fifoGroup_42_io_availability;
  wire                fifoGroup_43_io_push_ready;
  wire                fifoGroup_43_io_pop_valid;
  wire       [31:0]   fifoGroup_43_io_pop_payload;
  wire       [6:0]    fifoGroup_43_io_occupancy;
  wire       [6:0]    fifoGroup_43_io_availability;
  wire                fifoGroup_44_io_push_ready;
  wire                fifoGroup_44_io_pop_valid;
  wire       [31:0]   fifoGroup_44_io_pop_payload;
  wire       [6:0]    fifoGroup_44_io_occupancy;
  wire       [6:0]    fifoGroup_44_io_availability;
  wire                fifoGroup_45_io_push_ready;
  wire                fifoGroup_45_io_pop_valid;
  wire       [31:0]   fifoGroup_45_io_pop_payload;
  wire       [6:0]    fifoGroup_45_io_occupancy;
  wire       [6:0]    fifoGroup_45_io_availability;
  wire                fifoGroup_46_io_push_ready;
  wire                fifoGroup_46_io_pop_valid;
  wire       [31:0]   fifoGroup_46_io_pop_payload;
  wire       [6:0]    fifoGroup_46_io_occupancy;
  wire       [6:0]    fifoGroup_46_io_availability;
  wire                fifoGroup_47_io_push_ready;
  wire                fifoGroup_47_io_pop_valid;
  wire       [31:0]   fifoGroup_47_io_pop_payload;
  wire       [6:0]    fifoGroup_47_io_occupancy;
  wire       [6:0]    fifoGroup_47_io_availability;
  wire                fifoGroup_48_io_push_ready;
  wire                fifoGroup_48_io_pop_valid;
  wire       [31:0]   fifoGroup_48_io_pop_payload;
  wire       [6:0]    fifoGroup_48_io_occupancy;
  wire       [6:0]    fifoGroup_48_io_availability;
  wire                fifoGroup_49_io_push_ready;
  wire                fifoGroup_49_io_pop_valid;
  wire       [31:0]   fifoGroup_49_io_pop_payload;
  wire       [6:0]    fifoGroup_49_io_occupancy;
  wire       [6:0]    fifoGroup_49_io_availability;
  wire                fifoGroup_50_io_push_ready;
  wire                fifoGroup_50_io_pop_valid;
  wire       [31:0]   fifoGroup_50_io_pop_payload;
  wire       [6:0]    fifoGroup_50_io_occupancy;
  wire       [6:0]    fifoGroup_50_io_availability;
  wire                fifoGroup_51_io_push_ready;
  wire                fifoGroup_51_io_pop_valid;
  wire       [31:0]   fifoGroup_51_io_pop_payload;
  wire       [6:0]    fifoGroup_51_io_occupancy;
  wire       [6:0]    fifoGroup_51_io_availability;
  wire                fifoGroup_52_io_push_ready;
  wire                fifoGroup_52_io_pop_valid;
  wire       [31:0]   fifoGroup_52_io_pop_payload;
  wire       [6:0]    fifoGroup_52_io_occupancy;
  wire       [6:0]    fifoGroup_52_io_availability;
  wire                fifoGroup_53_io_push_ready;
  wire                fifoGroup_53_io_pop_valid;
  wire       [31:0]   fifoGroup_53_io_pop_payload;
  wire       [6:0]    fifoGroup_53_io_occupancy;
  wire       [6:0]    fifoGroup_53_io_availability;
  wire                fifoGroup_54_io_push_ready;
  wire                fifoGroup_54_io_pop_valid;
  wire       [31:0]   fifoGroup_54_io_pop_payload;
  wire       [6:0]    fifoGroup_54_io_occupancy;
  wire       [6:0]    fifoGroup_54_io_availability;
  wire                fifoGroup_55_io_push_ready;
  wire                fifoGroup_55_io_pop_valid;
  wire       [31:0]   fifoGroup_55_io_pop_payload;
  wire       [6:0]    fifoGroup_55_io_occupancy;
  wire       [6:0]    fifoGroup_55_io_availability;
  wire                fifoGroup_56_io_push_ready;
  wire                fifoGroup_56_io_pop_valid;
  wire       [31:0]   fifoGroup_56_io_pop_payload;
  wire       [6:0]    fifoGroup_56_io_occupancy;
  wire       [6:0]    fifoGroup_56_io_availability;
  wire                fifoGroup_57_io_push_ready;
  wire                fifoGroup_57_io_pop_valid;
  wire       [31:0]   fifoGroup_57_io_pop_payload;
  wire       [6:0]    fifoGroup_57_io_occupancy;
  wire       [6:0]    fifoGroup_57_io_availability;
  wire                fifoGroup_58_io_push_ready;
  wire                fifoGroup_58_io_pop_valid;
  wire       [31:0]   fifoGroup_58_io_pop_payload;
  wire       [6:0]    fifoGroup_58_io_occupancy;
  wire       [6:0]    fifoGroup_58_io_availability;
  wire                fifoGroup_59_io_push_ready;
  wire                fifoGroup_59_io_pop_valid;
  wire       [31:0]   fifoGroup_59_io_pop_payload;
  wire       [6:0]    fifoGroup_59_io_occupancy;
  wire       [6:0]    fifoGroup_59_io_availability;
  wire                fifoGroup_60_io_push_ready;
  wire                fifoGroup_60_io_pop_valid;
  wire       [31:0]   fifoGroup_60_io_pop_payload;
  wire       [6:0]    fifoGroup_60_io_occupancy;
  wire       [6:0]    fifoGroup_60_io_availability;
  wire                fifoGroup_61_io_push_ready;
  wire                fifoGroup_61_io_pop_valid;
  wire       [31:0]   fifoGroup_61_io_pop_payload;
  wire       [6:0]    fifoGroup_61_io_occupancy;
  wire       [6:0]    fifoGroup_61_io_availability;
  wire                fifoGroup_62_io_push_ready;
  wire                fifoGroup_62_io_pop_valid;
  wire       [31:0]   fifoGroup_62_io_pop_payload;
  wire       [6:0]    fifoGroup_62_io_occupancy;
  wire       [6:0]    fifoGroup_62_io_availability;
  wire                fifoGroup_63_io_push_ready;
  wire                fifoGroup_63_io_pop_valid;
  wire       [31:0]   fifoGroup_63_io_pop_payload;
  wire       [6:0]    fifoGroup_63_io_occupancy;
  wire       [6:0]    fifoGroup_63_io_availability;
  wire       [12:0]   _zz_handshakeTimes_0_valueNext;
  wire       [0:0]    _zz_handshakeTimes_0_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_1_valueNext;
  wire       [0:0]    _zz_handshakeTimes_1_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_2_valueNext;
  wire       [0:0]    _zz_handshakeTimes_2_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_3_valueNext;
  wire       [0:0]    _zz_handshakeTimes_3_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_4_valueNext;
  wire       [0:0]    _zz_handshakeTimes_4_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_5_valueNext;
  wire       [0:0]    _zz_handshakeTimes_5_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_6_valueNext;
  wire       [0:0]    _zz_handshakeTimes_6_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_7_valueNext;
  wire       [0:0]    _zz_handshakeTimes_7_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_0_valueNext;
  wire       [0:0]    _zz_outSliceNumb_0_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_1_valueNext;
  wire       [0:0]    _zz_outSliceNumb_1_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_2_valueNext;
  wire       [0:0]    _zz_outSliceNumb_2_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_3_valueNext;
  wire       [0:0]    _zz_outSliceNumb_3_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_4_valueNext;
  wire       [0:0]    _zz_outSliceNumb_4_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_5_valueNext;
  wire       [0:0]    _zz_outSliceNumb_5_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_6_valueNext;
  wire       [0:0]    _zz_outSliceNumb_6_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_7_valueNext;
  wire       [0:0]    _zz_outSliceNumb_7_valueNext_1;
  reg        [6:0]    _zz_when_ArraySlice_l211;
  wire       [6:0]    _zz_when_ArraySlice_l211_1;
  reg                 _zz_inputStreamArrayData_ready;
  reg        [6:0]    _zz_when_ArraySlice_l215;
  wire       [6:0]    _zz_when_ArraySlice_l215_1;
  wire       [5:0]    _zz_when_ArraySlice_l215_2;
  wire       [5:0]    _zz_when_ArraySlice_l215_3;
  wire       [0:0]    _zz_when_ArraySlice_l215_4;
  wire       [5:0]    _zz_when_ArraySlice_l216;
  wire       [5:0]    _zz_when_ArraySlice_l216_1;
  wire       [0:0]    _zz_when_ArraySlice_l216_2;
  wire       [5:0]    _zz_selectWriteFifo;
  wire       [0:0]    _zz_selectWriteFifo_1;
  wire       [5:0]    _zz_when_ArraySlice_l165;
  wire       [5:0]    _zz_when_ArraySlice_l165_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_2;
  wire       [6:0]    _zz_when_ArraySlice_l166;
  wire       [6:0]    _zz_when_ArraySlice_l166_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112;
  wire       [6:0]    _zz_when_ArraySlice_l113;
  wire       [6:0]    _zz_when_ArraySlice_l113_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_3;
  wire       [5:0]    _zz_when_ArraySlice_l118;
  wire       [6:0]    _zz_when_ArraySlice_l118_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_416;
  wire       [6:0]    _zz_when_ArraySlice_l173_417;
  wire       [6:0]    _zz_when_ArraySlice_l173_418;
  wire       [6:0]    _zz_when_ArraySlice_l173_419;
  wire       [5:0]    _zz_when_ArraySlice_l173_420;
  wire       [5:0]    _zz_when_ArraySlice_l173_421;
  wire       [2:0]    _zz_when_ArraySlice_l173_422;
  wire       [6:0]    _zz_when_ArraySlice_l173_423;
  wire       [5:0]    _zz_when_ArraySlice_l165_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l165_1_2;
  wire       [3:0]    _zz_when_ArraySlice_l165_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_1_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_1_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_1_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_1_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_1_4;
  wire       [6:0]    _zz_when_ArraySlice_l113_1_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_1_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_1_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_1_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l118_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l118_1_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_1_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_1_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_1_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_1_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_1_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_1_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_1_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_1_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l165_2_2;
  wire       [4:0]    _zz_when_ArraySlice_l165_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_2_4;
  wire       [4:0]    _zz_when_ArraySlice_l166_2_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_2_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_2_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_2_4;
  wire       [6:0]    _zz_when_ArraySlice_l113_2_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_2_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_2_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_2_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l118_2;
  wire       [6:0]    _zz_when_ArraySlice_l118_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_2_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_2_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_2_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_2_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_2_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_2_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_2_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_2_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_3;
  wire       [5:0]    _zz_when_ArraySlice_l165_3_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_3_4;
  wire       [4:0]    _zz_when_ArraySlice_l166_3_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_3_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_3_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_3_4;
  wire       [6:0]    _zz_when_ArraySlice_l113_3_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_3_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_3_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_3_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l118_3;
  wire       [6:0]    _zz_when_ArraySlice_l118_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_3_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_3_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_3_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_3_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_3_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_3_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_3_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_3_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_4;
  wire       [5:0]    _zz_when_ArraySlice_l165_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_4_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_4;
  wire       [6:0]    _zz_when_ArraySlice_l113_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_4_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_4_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l113_4_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_4_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_4_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_4;
  wire       [6:0]    _zz_when_ArraySlice_l118_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_4_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_4_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_4_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_4_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_4_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_4_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_5;
  wire       [5:0]    _zz_when_ArraySlice_l165_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_5_1;
  wire       [4:0]    _zz_when_ArraySlice_l166_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_5_4;
  wire       [5:0]    _zz_when_ArraySlice_l166_5_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_5;
  wire       [6:0]    _zz_when_ArraySlice_l113_5;
  wire       [6:0]    _zz_when_ArraySlice_l113_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_5_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_5_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_5_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_5_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_5;
  wire       [6:0]    _zz_when_ArraySlice_l118_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_5_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_5_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_5_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_5_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_5_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_5_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_5_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_6;
  wire       [5:0]    _zz_when_ArraySlice_l165_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_6;
  wire       [4:0]    _zz_when_ArraySlice_l166_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_6_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_6;
  wire       [6:0]    _zz_when_ArraySlice_l113_6;
  wire       [6:0]    _zz_when_ArraySlice_l113_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_6_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_6_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_6;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_6_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_6_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_6;
  wire       [6:0]    _zz_when_ArraySlice_l118_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_6_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_6_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_6_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_6_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_6_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_6_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_6_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_7;
  wire       [5:0]    _zz_when_ArraySlice_l165_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_7;
  wire       [3:0]    _zz_when_ArraySlice_l166_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_7_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_7;
  wire       [6:0]    _zz_when_ArraySlice_l113_7;
  wire       [6:0]    _zz_when_ArraySlice_l113_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_7_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_7_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_7;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_7_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_7_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_7;
  wire       [6:0]    _zz_when_ArraySlice_l118_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_7_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_7_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_7_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_7_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_7_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_7_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_7_8;
  wire       [5:0]    _zz_when_ArraySlice_l373;
  wire       [5:0]    _zz_when_ArraySlice_l373_1;
  wire       [2:0]    _zz_when_ArraySlice_l373_2;
  reg        [6:0]    _zz_when_ArraySlice_l374;
  wire       [5:0]    _zz_when_ArraySlice_l374_1;
  wire       [5:0]    _zz_when_ArraySlice_l374_2;
  wire       [2:0]    _zz_when_ArraySlice_l374_3;
  wire       [5:0]    _zz__zz_outputStreamArrayData_0_valid;
  wire       [2:0]    _zz__zz_outputStreamArrayData_0_valid_1;
  reg                 _zz_outputStreamArrayData_0_valid_2;
  reg        [31:0]   _zz_outputStreamArrayData_0_payload;
  wire       [6:0]    _zz_when_ArraySlice_l380;
  wire       [0:0]    _zz_when_ArraySlice_l380_1;
  reg        [6:0]    _zz_when_ArraySlice_l380_2;
  wire       [5:0]    _zz_when_ArraySlice_l380_3;
  wire       [5:0]    _zz_when_ArraySlice_l380_4;
  wire       [2:0]    _zz_when_ArraySlice_l380_5;
  wire       [12:0]   _zz_when_ArraySlice_l381;
  wire       [5:0]    _zz_when_ArraySlice_l381_1;
  wire       [5:0]    _zz_when_ArraySlice_l381_2;
  wire       [5:0]    _zz_when_ArraySlice_l381_3;
  wire       [0:0]    _zz_when_ArraySlice_l381_4;
  wire       [5:0]    _zz_selectReadFifo_0;
  wire       [5:0]    _zz_selectReadFifo_0_1;
  wire       [5:0]    _zz_selectReadFifo_0_2;
  wire       [0:0]    _zz_selectReadFifo_0_3;
  wire       [5:0]    _zz_selectReadFifo_0_4;
  wire       [0:0]    _zz_selectReadFifo_0_5;
  wire       [12:0]   _zz_when_ArraySlice_l384;
  wire       [12:0]   _zz_when_ArraySlice_l384_1;
  wire       [12:0]   _zz_when_ArraySlice_l384_2;
  wire       [0:0]    _zz_when_ArraySlice_l384_3;
  reg        [6:0]    _zz_when_ArraySlice_l389;
  wire       [5:0]    _zz_when_ArraySlice_l389_1;
  wire       [5:0]    _zz_when_ArraySlice_l389_2;
  wire       [2:0]    _zz_when_ArraySlice_l389_3;
  wire       [6:0]    _zz_when_ArraySlice_l389_4;
  wire       [0:0]    _zz_when_ArraySlice_l389_5;
  wire       [12:0]   _zz_when_ArraySlice_l390;
  wire       [5:0]    _zz_when_ArraySlice_l390_1;
  wire       [5:0]    _zz_when_ArraySlice_l390_2;
  wire       [5:0]    _zz_when_ArraySlice_l390_3;
  wire       [0:0]    _zz_when_ArraySlice_l390_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94;
  wire       [6:0]    _zz_when_ArraySlice_l95;
  wire       [6:0]    _zz_when_ArraySlice_l95_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_3;
  wire       [5:0]    _zz_when_ArraySlice_l99;
  wire       [6:0]    _zz_when_ArraySlice_l99_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_8;
  wire       [6:0]    _zz_when_ArraySlice_l392_9;
  wire       [0:0]    _zz_when_ArraySlice_l392_10;
  wire       [6:0]    _zz_when_ArraySlice_l392_11;
  wire       [5:0]    _zz_selectReadFifo_0_6;
  wire       [5:0]    _zz_selectReadFifo_0_7;
  wire       [5:0]    _zz_selectReadFifo_0_8;
  wire       [0:0]    _zz_selectReadFifo_0_9;
  wire       [5:0]    _zz_selectReadFifo_0_10;
  wire       [5:0]    _zz_selectReadFifo_0_11;
  wire       [5:0]    _zz_selectReadFifo_0_12;
  wire       [0:0]    _zz_selectReadFifo_0_13;
  wire       [5:0]    _zz_when_ArraySlice_l165_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_8_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_8_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_8;
  wire       [6:0]    _zz_when_ArraySlice_l166_8_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_8_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_8_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_8_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_8_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_8;
  wire       [6:0]    _zz_when_ArraySlice_l113_8;
  wire       [6:0]    _zz_when_ArraySlice_l113_8_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_8_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_8_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_8_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_8;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_8_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_8_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_8_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_8;
  wire       [6:0]    _zz_when_ArraySlice_l118_8_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_8_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_8_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_8_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_8_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_8_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_8_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_8_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_8_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_9_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_9_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_9;
  wire       [5:0]    _zz_when_ArraySlice_l166_9_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_9_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_9_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_9_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_9;
  wire       [6:0]    _zz_when_ArraySlice_l113_9;
  wire       [6:0]    _zz_when_ArraySlice_l113_9_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_9_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_9_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_9_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_9;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_9_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_9_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_9_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_9;
  wire       [6:0]    _zz_when_ArraySlice_l118_9_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_9_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_9_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_9_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_9_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_9_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_9_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_9_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_9_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_9_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_10;
  wire       [5:0]    _zz_when_ArraySlice_l165_10_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_10_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_10;
  wire       [5:0]    _zz_when_ArraySlice_l166_10_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_10_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_10_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_10_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_10;
  wire       [6:0]    _zz_when_ArraySlice_l113_10;
  wire       [6:0]    _zz_when_ArraySlice_l113_10_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_10_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_10_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_10_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_10;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_10_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_10_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_10_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_10;
  wire       [6:0]    _zz_when_ArraySlice_l118_10_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_10_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_10_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_10_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_10_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_10_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_10_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_10_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_10_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_10_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_11;
  wire       [5:0]    _zz_when_ArraySlice_l165_11_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_11_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_11;
  wire       [5:0]    _zz_when_ArraySlice_l166_11_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_11_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_11_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_11_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_11;
  wire       [6:0]    _zz_when_ArraySlice_l113_11;
  wire       [6:0]    _zz_when_ArraySlice_l113_11_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_11_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_11_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_11_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_11;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_11_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_11_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_11_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_11;
  wire       [6:0]    _zz_when_ArraySlice_l118_11_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_11_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_11_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_11_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_11_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_11_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_11_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_11_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_11_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_11_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_12;
  wire       [5:0]    _zz_when_ArraySlice_l165_12_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_12;
  wire       [5:0]    _zz_when_ArraySlice_l166_12_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_12_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_12_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_12;
  wire       [6:0]    _zz_when_ArraySlice_l113_12;
  wire       [6:0]    _zz_when_ArraySlice_l113_12_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_12_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_12_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_12_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_12;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_12_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_12_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_12_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_12;
  wire       [6:0]    _zz_when_ArraySlice_l118_12_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_12_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_12_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_12_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_12_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_12_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_12_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_12_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_12_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_13;
  wire       [5:0]    _zz_when_ArraySlice_l165_13_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_13;
  wire       [4:0]    _zz_when_ArraySlice_l166_13_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_13_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_13_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_13_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_13;
  wire       [6:0]    _zz_when_ArraySlice_l113_13;
  wire       [6:0]    _zz_when_ArraySlice_l113_13_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_13_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_13_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_13_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_13;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_13_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_13_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_13_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_13;
  wire       [6:0]    _zz_when_ArraySlice_l118_13_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_13_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_13_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_13_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_13_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_13_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_13_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_13_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_13_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_14;
  wire       [5:0]    _zz_when_ArraySlice_l165_14_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_14;
  wire       [4:0]    _zz_when_ArraySlice_l166_14_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_14_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_14_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_14_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_14;
  wire       [6:0]    _zz_when_ArraySlice_l113_14;
  wire       [6:0]    _zz_when_ArraySlice_l113_14_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_14_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_14_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_14_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_14;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_14_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_14_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_14_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_14;
  wire       [6:0]    _zz_when_ArraySlice_l118_14_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_14_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_14_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_14_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_14_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_14_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_14_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_14_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_14_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_15;
  wire       [5:0]    _zz_when_ArraySlice_l165_15_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_15;
  wire       [3:0]    _zz_when_ArraySlice_l166_15_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_15_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_15_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_15_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_15;
  wire       [6:0]    _zz_when_ArraySlice_l113_15;
  wire       [6:0]    _zz_when_ArraySlice_l113_15_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_15_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_15_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_15_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_15;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_15_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_15_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_15_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_15;
  wire       [6:0]    _zz_when_ArraySlice_l118_15_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_15_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_15_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_15_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_15_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_15_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_15_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_15_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_15_8;
  wire                _zz_when_ArraySlice_l398;
  wire                _zz_when_ArraySlice_l398_1;
  wire                _zz_when_ArraySlice_l398_2;
  wire                _zz_when_ArraySlice_l398_3;
  wire                _zz_when_ArraySlice_l398_4;
  wire                _zz_when_ArraySlice_l398_5;
  wire                _zz_when_ArraySlice_l398_6;
  wire                _zz_when_ArraySlice_l398_7;
  wire                _zz_when_ArraySlice_l398_8;
  wire                _zz_when_ArraySlice_l398_9;
  wire       [5:0]    _zz_when_ArraySlice_l401;
  wire       [5:0]    _zz_when_ArraySlice_l401_1;
  wire       [5:0]    _zz_when_ArraySlice_l401_2;
  wire       [5:0]    _zz_when_ArraySlice_l401_3;
  wire       [5:0]    _zz_when_ArraySlice_l401_4;
  wire       [0:0]    _zz_when_ArraySlice_l401_5;
  wire       [5:0]    _zz_when_ArraySlice_l401_6;
  wire       [2:0]    _zz_when_ArraySlice_l401_7;
  wire       [5:0]    _zz_selectReadFifo_0_14;
  wire       [0:0]    _zz_selectReadFifo_0_15;
  wire       [12:0]   _zz_when_ArraySlice_l405;
  wire       [12:0]   _zz_when_ArraySlice_l405_1;
  wire       [12:0]   _zz_when_ArraySlice_l405_2;
  wire       [0:0]    _zz_when_ArraySlice_l405_3;
  reg        [6:0]    _zz_when_ArraySlice_l409;
  wire       [5:0]    _zz_when_ArraySlice_l409_1;
  wire       [5:0]    _zz_when_ArraySlice_l409_2;
  wire       [2:0]    _zz_when_ArraySlice_l409_3;
  wire       [12:0]   _zz_when_ArraySlice_l410;
  wire       [5:0]    _zz_when_ArraySlice_l410_1;
  wire       [5:0]    _zz_when_ArraySlice_l410_2;
  wire       [5:0]    _zz_when_ArraySlice_l410_3;
  wire       [0:0]    _zz_when_ArraySlice_l410_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_1_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_1_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_1_4;
  wire       [6:0]    _zz_when_ArraySlice_l95_1_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l99_1_2;
  wire       [6:0]    _zz_when_ArraySlice_l412_8;
  wire       [6:0]    _zz_when_ArraySlice_l412_9;
  wire       [0:0]    _zz_when_ArraySlice_l412_10;
  wire       [6:0]    _zz_when_ArraySlice_l412_11;
  wire       [5:0]    _zz_selectReadFifo_0_16;
  wire       [5:0]    _zz_selectReadFifo_0_17;
  wire       [5:0]    _zz_selectReadFifo_0_18;
  wire       [0:0]    _zz_selectReadFifo_0_19;
  wire       [5:0]    _zz_selectReadFifo_0_20;
  wire       [5:0]    _zz_selectReadFifo_0_21;
  wire       [5:0]    _zz_selectReadFifo_0_22;
  wire       [0:0]    _zz_selectReadFifo_0_23;
  wire       [5:0]    _zz_when_ArraySlice_l165_16;
  wire       [5:0]    _zz_when_ArraySlice_l165_16_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_16_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_16;
  wire       [6:0]    _zz_when_ArraySlice_l166_16_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_16_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_16_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_16_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_16_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_16;
  wire       [6:0]    _zz_when_ArraySlice_l113_16;
  wire       [6:0]    _zz_when_ArraySlice_l113_16_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_16_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_16_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_16_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_16;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_16_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_16_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_16_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_16;
  wire       [6:0]    _zz_when_ArraySlice_l118_16_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_16_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_16_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_16_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_16_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_16_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_16_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_16_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_16_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_17;
  wire       [5:0]    _zz_when_ArraySlice_l165_17_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_17_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_17;
  wire       [5:0]    _zz_when_ArraySlice_l166_17_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_17_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_17_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_17_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_17;
  wire       [6:0]    _zz_when_ArraySlice_l113_17;
  wire       [6:0]    _zz_when_ArraySlice_l113_17_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_17_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_17_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_17_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_17;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_17_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_17_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_17_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_17;
  wire       [6:0]    _zz_when_ArraySlice_l118_17_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_17_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_17_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_17_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_17_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_17_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_17_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_17_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_17_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_17_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_18;
  wire       [5:0]    _zz_when_ArraySlice_l165_18_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_18_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_18;
  wire       [5:0]    _zz_when_ArraySlice_l166_18_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_18_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_18_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_18_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_18;
  wire       [6:0]    _zz_when_ArraySlice_l113_18;
  wire       [6:0]    _zz_when_ArraySlice_l113_18_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_18_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_18_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_18_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_18;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_18_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_18_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_18_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_18;
  wire       [6:0]    _zz_when_ArraySlice_l118_18_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_18_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_18_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_18_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_18_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_18_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_18_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_18_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_18_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_18_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_19;
  wire       [5:0]    _zz_when_ArraySlice_l165_19_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_19_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_19;
  wire       [5:0]    _zz_when_ArraySlice_l166_19_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_19_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_19_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_19_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_19;
  wire       [6:0]    _zz_when_ArraySlice_l113_19;
  wire       [6:0]    _zz_when_ArraySlice_l113_19_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_19_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_19_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_19_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_19;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_19_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_19_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_19_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_19;
  wire       [6:0]    _zz_when_ArraySlice_l118_19_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_19_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_19_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_19_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_19_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_19_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_19_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_19_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_19_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_19_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_20;
  wire       [5:0]    _zz_when_ArraySlice_l165_20_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_20;
  wire       [5:0]    _zz_when_ArraySlice_l166_20_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_20_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_20_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_20;
  wire       [6:0]    _zz_when_ArraySlice_l113_20;
  wire       [6:0]    _zz_when_ArraySlice_l113_20_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_20_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_20_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_20_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_20;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_20_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_20_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_20_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_20;
  wire       [6:0]    _zz_when_ArraySlice_l118_20_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_20_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_20_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_20_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_20_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_20_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_20_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_20_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_20_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_21;
  wire       [5:0]    _zz_when_ArraySlice_l165_21_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_21;
  wire       [4:0]    _zz_when_ArraySlice_l166_21_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_21_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_21_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_21_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_21;
  wire       [6:0]    _zz_when_ArraySlice_l113_21;
  wire       [6:0]    _zz_when_ArraySlice_l113_21_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_21_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_21_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_21_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_21;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_21_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_21_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_21_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_21;
  wire       [6:0]    _zz_when_ArraySlice_l118_21_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_21_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_21_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_21_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_21_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_21_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_21_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_21_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_21_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_22;
  wire       [5:0]    _zz_when_ArraySlice_l165_22_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_22;
  wire       [4:0]    _zz_when_ArraySlice_l166_22_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_22_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_22_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_22_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_22;
  wire       [6:0]    _zz_when_ArraySlice_l113_22;
  wire       [6:0]    _zz_when_ArraySlice_l113_22_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_22_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_22_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_22_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_22;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_22_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_22_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_22_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_22;
  wire       [6:0]    _zz_when_ArraySlice_l118_22_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_22_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_22_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_22_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_22_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_22_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_22_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_22_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_22_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_23;
  wire       [5:0]    _zz_when_ArraySlice_l165_23_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_23;
  wire       [3:0]    _zz_when_ArraySlice_l166_23_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_23_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_23_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_23_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_23;
  wire       [6:0]    _zz_when_ArraySlice_l113_23;
  wire       [6:0]    _zz_when_ArraySlice_l113_23_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_23_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_23_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_23_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_23;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_23_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_23_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_23_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_23;
  wire       [6:0]    _zz_when_ArraySlice_l118_23_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_23_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_23_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_23_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_23_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_23_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_23_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_23_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_23_8;
  wire                _zz_when_ArraySlice_l418;
  wire                _zz_when_ArraySlice_l418_1;
  wire                _zz_when_ArraySlice_l418_2;
  wire                _zz_when_ArraySlice_l418_3;
  wire                _zz_when_ArraySlice_l418_4;
  wire                _zz_when_ArraySlice_l418_5;
  wire       [5:0]    _zz_when_ArraySlice_l421;
  wire       [5:0]    _zz_when_ArraySlice_l421_1;
  wire       [5:0]    _zz_when_ArraySlice_l421_2;
  wire       [5:0]    _zz_when_ArraySlice_l421_3;
  wire       [5:0]    _zz_when_ArraySlice_l421_4;
  wire       [0:0]    _zz_when_ArraySlice_l421_5;
  wire       [5:0]    _zz_when_ArraySlice_l421_6;
  wire       [2:0]    _zz_when_ArraySlice_l421_7;
  wire       [5:0]    _zz_selectReadFifo_0_24;
  wire       [0:0]    _zz_selectReadFifo_0_25;
  wire       [12:0]   _zz_when_ArraySlice_l425;
  wire       [12:0]   _zz_when_ArraySlice_l425_1;
  wire       [12:0]   _zz_when_ArraySlice_l425_2;
  wire       [0:0]    _zz_when_ArraySlice_l425_3;
  wire       [12:0]   _zz_when_ArraySlice_l436;
  wire       [5:0]    _zz_when_ArraySlice_l436_1;
  wire       [5:0]    _zz_when_ArraySlice_l436_2;
  wire       [5:0]    _zz_when_ArraySlice_l436_3;
  wire       [0:0]    _zz_when_ArraySlice_l436_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_2_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_2_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_2_4;
  wire       [6:0]    _zz_when_ArraySlice_l95_2_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_2;
  wire       [6:0]    _zz_when_ArraySlice_l99_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_8;
  wire       [6:0]    _zz_when_ArraySlice_l437_9;
  wire       [0:0]    _zz_when_ArraySlice_l437_10;
  wire       [6:0]    _zz_when_ArraySlice_l437_11;
  wire       [5:0]    _zz_selectReadFifo_0_26;
  wire       [5:0]    _zz_selectReadFifo_0_27;
  wire       [5:0]    _zz_selectReadFifo_0_28;
  wire       [0:0]    _zz_selectReadFifo_0_29;
  wire       [5:0]    _zz_when_ArraySlice_l165_24;
  wire       [5:0]    _zz_when_ArraySlice_l165_24_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_24_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_24;
  wire       [6:0]    _zz_when_ArraySlice_l166_24_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_24_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_24_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_24_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_24_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_24;
  wire       [6:0]    _zz_when_ArraySlice_l113_24;
  wire       [6:0]    _zz_when_ArraySlice_l113_24_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_24_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_24_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_24_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_24;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_24_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_24_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_24_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_24;
  wire       [6:0]    _zz_when_ArraySlice_l118_24_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_24_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_24_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_24_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_24_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_24_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_24_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_24_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_24_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_25;
  wire       [5:0]    _zz_when_ArraySlice_l165_25_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_25_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_25;
  wire       [5:0]    _zz_when_ArraySlice_l166_25_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_25_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_25_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_25_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_25;
  wire       [6:0]    _zz_when_ArraySlice_l113_25;
  wire       [6:0]    _zz_when_ArraySlice_l113_25_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_25_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_25_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_25_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_25;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_25_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_25_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_25_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_25;
  wire       [6:0]    _zz_when_ArraySlice_l118_25_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_25_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_25_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_25_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_25_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_25_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_25_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_25_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_25_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_25_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_26;
  wire       [5:0]    _zz_when_ArraySlice_l165_26_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_26_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_26;
  wire       [5:0]    _zz_when_ArraySlice_l166_26_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_26_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_26_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_26_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_26;
  wire       [6:0]    _zz_when_ArraySlice_l113_26;
  wire       [6:0]    _zz_when_ArraySlice_l113_26_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_26_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_26_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_26_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_26;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_26_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_26_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_26_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_26;
  wire       [6:0]    _zz_when_ArraySlice_l118_26_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_26_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_26_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_26_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_26_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_26_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_26_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_26_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_26_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_26_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_27;
  wire       [5:0]    _zz_when_ArraySlice_l165_27_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_27_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_27;
  wire       [5:0]    _zz_when_ArraySlice_l166_27_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_27_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_27_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_27_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_27;
  wire       [6:0]    _zz_when_ArraySlice_l113_27;
  wire       [6:0]    _zz_when_ArraySlice_l113_27_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_27_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_27_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_27_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_27;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_27_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_27_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_27_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_27;
  wire       [6:0]    _zz_when_ArraySlice_l118_27_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_27_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_27_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_27_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_27_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_27_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_27_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_27_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_27_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_27_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_28;
  wire       [5:0]    _zz_when_ArraySlice_l165_28_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_28;
  wire       [5:0]    _zz_when_ArraySlice_l166_28_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_28_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_28_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_28;
  wire       [6:0]    _zz_when_ArraySlice_l113_28;
  wire       [6:0]    _zz_when_ArraySlice_l113_28_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_28_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_28_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_28_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_28;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_28_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_28_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_28_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_28;
  wire       [6:0]    _zz_when_ArraySlice_l118_28_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_28_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_28_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_28_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_28_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_28_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_28_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_28_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_28_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_29;
  wire       [5:0]    _zz_when_ArraySlice_l165_29_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_29;
  wire       [4:0]    _zz_when_ArraySlice_l166_29_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_29_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_29_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_29_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_29;
  wire       [6:0]    _zz_when_ArraySlice_l113_29;
  wire       [6:0]    _zz_when_ArraySlice_l113_29_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_29_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_29_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_29_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_29;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_29_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_29_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_29_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_29;
  wire       [6:0]    _zz_when_ArraySlice_l118_29_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_29_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_29_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_29_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_29_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_29_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_29_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_29_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_29_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_30;
  wire       [5:0]    _zz_when_ArraySlice_l165_30_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_30;
  wire       [4:0]    _zz_when_ArraySlice_l166_30_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_30_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_30_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_30_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_30;
  wire       [6:0]    _zz_when_ArraySlice_l113_30;
  wire       [6:0]    _zz_when_ArraySlice_l113_30_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_30_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_30_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_30_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_30;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_30_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_30_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_30_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_30;
  wire       [6:0]    _zz_when_ArraySlice_l118_30_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_30_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_30_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_30_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_30_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_30_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_30_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_30_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_30_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_31;
  wire       [5:0]    _zz_when_ArraySlice_l165_31_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_31;
  wire       [3:0]    _zz_when_ArraySlice_l166_31_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_31_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_31_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_31_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_31;
  wire       [6:0]    _zz_when_ArraySlice_l113_31;
  wire       [6:0]    _zz_when_ArraySlice_l113_31_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_31_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_31_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_31_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_31;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_31_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_31_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_31_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_31;
  wire       [6:0]    _zz_when_ArraySlice_l118_31_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_31_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_31_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_31_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_31_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_31_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_31_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_31_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_31_8;
  wire                _zz_when_ArraySlice_l444;
  wire                _zz_when_ArraySlice_l444_1;
  wire                _zz_when_ArraySlice_l444_2;
  wire                _zz_when_ArraySlice_l444_3;
  wire                _zz_when_ArraySlice_l444_4;
  wire                _zz_when_ArraySlice_l444_5;
  wire       [5:0]    _zz_selectReadFifo_0_30;
  wire       [0:0]    _zz_selectReadFifo_0_31;
  wire       [12:0]   _zz_when_ArraySlice_l448;
  wire       [12:0]   _zz_when_ArraySlice_l448_1;
  wire       [12:0]   _zz_when_ArraySlice_l448_2;
  wire       [0:0]    _zz_when_ArraySlice_l448_3;
  wire       [5:0]    _zz_when_ArraySlice_l434;
  wire       [5:0]    _zz_when_ArraySlice_l434_1;
  wire       [2:0]    _zz_when_ArraySlice_l434_2;
  wire       [12:0]   _zz_when_ArraySlice_l455;
  wire       [5:0]    _zz_when_ArraySlice_l455_1;
  wire       [5:0]    _zz_when_ArraySlice_l455_2;
  wire       [5:0]    _zz_when_ArraySlice_l455_3;
  wire       [0:0]    _zz_when_ArraySlice_l455_4;
  wire       [5:0]    _zz_when_ArraySlice_l373_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l373_1_2;
  wire       [3:0]    _zz_when_ArraySlice_l373_1_3;
  reg        [6:0]    _zz_when_ArraySlice_l374_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l374_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l374_1_3;
  wire       [3:0]    _zz_when_ArraySlice_l374_1_4;
  wire       [5:0]    _zz__zz_outputStreamArrayData_1_valid;
  wire       [3:0]    _zz__zz_outputStreamArrayData_1_valid_1;
  reg                 _zz_outputStreamArrayData_1_valid_2;
  reg        [31:0]   _zz_outputStreamArrayData_1_payload;
  wire       [6:0]    _zz_when_ArraySlice_l380_1_1;
  wire       [0:0]    _zz_when_ArraySlice_l380_1_2;
  reg        [6:0]    _zz_when_ArraySlice_l380_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l380_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l380_1_5;
  wire       [3:0]    _zz_when_ArraySlice_l380_1_6;
  wire       [12:0]   _zz_when_ArraySlice_l381_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l381_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l381_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l381_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l381_1_5;
  wire       [5:0]    _zz_selectReadFifo_1;
  wire       [5:0]    _zz_selectReadFifo_1_1;
  wire       [5:0]    _zz_selectReadFifo_1_2;
  wire       [0:0]    _zz_selectReadFifo_1_3;
  wire       [5:0]    _zz_selectReadFifo_1_4;
  wire       [0:0]    _zz_selectReadFifo_1_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l384_1_2;
  wire       [12:0]   _zz_when_ArraySlice_l384_1_3;
  wire       [0:0]    _zz_when_ArraySlice_l384_1_4;
  reg        [6:0]    _zz_when_ArraySlice_l389_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l389_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l389_1_3;
  wire       [3:0]    _zz_when_ArraySlice_l389_1_4;
  wire       [6:0]    _zz_when_ArraySlice_l389_1_5;
  wire       [0:0]    _zz_when_ArraySlice_l389_1_6;
  wire       [12:0]   _zz_when_ArraySlice_l390_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l390_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l390_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l390_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l390_1_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_3_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_3_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_3_4;
  wire       [6:0]    _zz_when_ArraySlice_l95_3_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_1_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_1_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_1_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_3;
  wire       [6:0]    _zz_when_ArraySlice_l99_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_1_2;
  wire       [0:0]    _zz_when_ArraySlice_l392_1_3;
  wire       [6:0]    _zz_when_ArraySlice_l392_1_4;
  wire       [5:0]    _zz_selectReadFifo_1_6;
  wire       [5:0]    _zz_selectReadFifo_1_7;
  wire       [5:0]    _zz_selectReadFifo_1_8;
  wire       [0:0]    _zz_selectReadFifo_1_9;
  wire       [5:0]    _zz_selectReadFifo_1_10;
  wire       [5:0]    _zz_selectReadFifo_1_11;
  wire       [5:0]    _zz_selectReadFifo_1_12;
  wire       [0:0]    _zz_selectReadFifo_1_13;
  wire       [5:0]    _zz_when_ArraySlice_l165_32;
  wire       [5:0]    _zz_when_ArraySlice_l165_32_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_32_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_32;
  wire       [6:0]    _zz_when_ArraySlice_l166_32_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_32_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_32_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_32_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_32_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_32;
  wire       [6:0]    _zz_when_ArraySlice_l113_32;
  wire       [6:0]    _zz_when_ArraySlice_l113_32_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_32_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_32_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_32_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_32;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_32_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_32_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_32_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_32;
  wire       [6:0]    _zz_when_ArraySlice_l118_32_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_32_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_32_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_32_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_32_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_32_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_32_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_32_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_32_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_33;
  wire       [5:0]    _zz_when_ArraySlice_l165_33_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_33_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_33;
  wire       [5:0]    _zz_when_ArraySlice_l166_33_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_33_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_33_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_33_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_33;
  wire       [6:0]    _zz_when_ArraySlice_l113_33;
  wire       [6:0]    _zz_when_ArraySlice_l113_33_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_33_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_33_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_33_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_33;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_33_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_33_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_33_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_33;
  wire       [6:0]    _zz_when_ArraySlice_l118_33_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_33_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_33_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_33_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_33_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_33_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_33_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_33_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_33_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_33_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_34;
  wire       [5:0]    _zz_when_ArraySlice_l165_34_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_34_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_34;
  wire       [5:0]    _zz_when_ArraySlice_l166_34_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_34_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_34_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_34_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_34;
  wire       [6:0]    _zz_when_ArraySlice_l113_34;
  wire       [6:0]    _zz_when_ArraySlice_l113_34_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_34_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_34_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_34_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_34;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_34_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_34_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_34_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_34;
  wire       [6:0]    _zz_when_ArraySlice_l118_34_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_34_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_34_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_34_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_34_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_34_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_34_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_34_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_34_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_34_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_35;
  wire       [5:0]    _zz_when_ArraySlice_l165_35_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_35_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_35;
  wire       [5:0]    _zz_when_ArraySlice_l166_35_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_35_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_35_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_35_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_35;
  wire       [6:0]    _zz_when_ArraySlice_l113_35;
  wire       [6:0]    _zz_when_ArraySlice_l113_35_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_35_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_35_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_35_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_35;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_35_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_35_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_35_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_35;
  wire       [6:0]    _zz_when_ArraySlice_l118_35_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_35_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_35_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_35_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_35_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_35_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_35_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_35_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_35_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_35_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_36;
  wire       [5:0]    _zz_when_ArraySlice_l165_36_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_36;
  wire       [5:0]    _zz_when_ArraySlice_l166_36_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_36_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_36_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_36;
  wire       [6:0]    _zz_when_ArraySlice_l113_36;
  wire       [6:0]    _zz_when_ArraySlice_l113_36_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_36_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_36_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_36_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_36;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_36_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_36_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_36_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_36;
  wire       [6:0]    _zz_when_ArraySlice_l118_36_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_36_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_36_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_36_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_36_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_36_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_36_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_36_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_36_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_37;
  wire       [5:0]    _zz_when_ArraySlice_l165_37_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_37;
  wire       [4:0]    _zz_when_ArraySlice_l166_37_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_37_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_37_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_37_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_37;
  wire       [6:0]    _zz_when_ArraySlice_l113_37;
  wire       [6:0]    _zz_when_ArraySlice_l113_37_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_37_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_37_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_37_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_37;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_37_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_37_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_37_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_37;
  wire       [6:0]    _zz_when_ArraySlice_l118_37_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_37_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_37_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_37_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_37_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_37_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_37_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_37_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_37_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_38;
  wire       [5:0]    _zz_when_ArraySlice_l165_38_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_38;
  wire       [4:0]    _zz_when_ArraySlice_l166_38_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_38_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_38_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_38_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_38;
  wire       [6:0]    _zz_when_ArraySlice_l113_38;
  wire       [6:0]    _zz_when_ArraySlice_l113_38_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_38_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_38_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_38_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_38;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_38_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_38_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_38_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_38;
  wire       [6:0]    _zz_when_ArraySlice_l118_38_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_38_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_38_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_38_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_38_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_38_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_38_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_38_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_38_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_39;
  wire       [5:0]    _zz_when_ArraySlice_l165_39_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_39;
  wire       [3:0]    _zz_when_ArraySlice_l166_39_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_39_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_39_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_39_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_39;
  wire       [6:0]    _zz_when_ArraySlice_l113_39;
  wire       [6:0]    _zz_when_ArraySlice_l113_39_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_39_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_39_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_39_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_39;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_39_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_39_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_39_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_39;
  wire       [6:0]    _zz_when_ArraySlice_l118_39_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_39_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_39_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_39_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_39_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_39_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_39_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_39_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_39_8;
  wire                _zz_when_ArraySlice_l398_1_1;
  wire                _zz_when_ArraySlice_l398_1_2;
  wire                _zz_when_ArraySlice_l398_1_3;
  wire                _zz_when_ArraySlice_l398_1_4;
  wire                _zz_when_ArraySlice_l398_1_5;
  wire                _zz_when_ArraySlice_l398_1_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l401_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l401_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l401_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l401_1_5;
  wire       [0:0]    _zz_when_ArraySlice_l401_1_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_1_7;
  wire       [3:0]    _zz_when_ArraySlice_l401_1_8;
  wire       [5:0]    _zz_selectReadFifo_1_14;
  wire       [0:0]    _zz_selectReadFifo_1_15;
  wire       [12:0]   _zz_when_ArraySlice_l405_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l405_1_2;
  wire       [12:0]   _zz_when_ArraySlice_l405_1_3;
  wire       [0:0]    _zz_when_ArraySlice_l405_1_4;
  reg        [6:0]    _zz_when_ArraySlice_l409_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l409_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l409_1_3;
  wire       [3:0]    _zz_when_ArraySlice_l409_1_4;
  wire       [12:0]   _zz_when_ArraySlice_l410_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l410_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l410_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l410_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l410_1_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_4;
  wire       [6:0]    _zz_when_ArraySlice_l95_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_4_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_4_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l95_4_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_1_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_1_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_1_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_4;
  wire       [6:0]    _zz_when_ArraySlice_l99_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_1_2;
  wire       [0:0]    _zz_when_ArraySlice_l412_1_3;
  wire       [6:0]    _zz_when_ArraySlice_l412_1_4;
  wire       [5:0]    _zz_selectReadFifo_1_16;
  wire       [5:0]    _zz_selectReadFifo_1_17;
  wire       [5:0]    _zz_selectReadFifo_1_18;
  wire       [0:0]    _zz_selectReadFifo_1_19;
  wire       [5:0]    _zz_selectReadFifo_1_20;
  wire       [5:0]    _zz_selectReadFifo_1_21;
  wire       [5:0]    _zz_selectReadFifo_1_22;
  wire       [0:0]    _zz_selectReadFifo_1_23;
  wire       [5:0]    _zz_when_ArraySlice_l165_40;
  wire       [5:0]    _zz_when_ArraySlice_l165_40_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_40_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_40;
  wire       [6:0]    _zz_when_ArraySlice_l166_40_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_40_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_40_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_40_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_40_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_40;
  wire       [6:0]    _zz_when_ArraySlice_l113_40;
  wire       [6:0]    _zz_when_ArraySlice_l113_40_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_40_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_40_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_40_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_40;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_40_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_40_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_40_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_40;
  wire       [6:0]    _zz_when_ArraySlice_l118_40_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_40_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_40_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_40_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_40_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_40_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_40_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_40_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_40_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_41;
  wire       [5:0]    _zz_when_ArraySlice_l165_41_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_41_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_41;
  wire       [5:0]    _zz_when_ArraySlice_l166_41_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_41_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_41_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_41_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_41;
  wire       [6:0]    _zz_when_ArraySlice_l113_41;
  wire       [6:0]    _zz_when_ArraySlice_l113_41_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_41_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_41_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_41_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_41;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_41_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_41_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_41_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_41;
  wire       [6:0]    _zz_when_ArraySlice_l118_41_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_41_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_41_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_41_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_41_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_41_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_41_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_41_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_41_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_41_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_42;
  wire       [5:0]    _zz_when_ArraySlice_l165_42_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_42_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_42;
  wire       [5:0]    _zz_when_ArraySlice_l166_42_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_42_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_42_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_42_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_42;
  wire       [6:0]    _zz_when_ArraySlice_l113_42;
  wire       [6:0]    _zz_when_ArraySlice_l113_42_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_42_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_42_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_42_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_42;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_42_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_42_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_42_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_42;
  wire       [6:0]    _zz_when_ArraySlice_l118_42_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_42_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_42_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_42_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_42_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_42_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_42_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_42_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_42_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_42_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_43;
  wire       [5:0]    _zz_when_ArraySlice_l165_43_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_43_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_43;
  wire       [5:0]    _zz_when_ArraySlice_l166_43_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_43_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_43_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_43_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_43;
  wire       [6:0]    _zz_when_ArraySlice_l113_43;
  wire       [6:0]    _zz_when_ArraySlice_l113_43_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_43_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_43_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_43_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_43;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_43_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_43_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_43_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_43;
  wire       [6:0]    _zz_when_ArraySlice_l118_43_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_43_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_43_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_43_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_43_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_43_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_43_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_43_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_43_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_43_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_44;
  wire       [5:0]    _zz_when_ArraySlice_l165_44_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_44;
  wire       [5:0]    _zz_when_ArraySlice_l166_44_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_44_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_44_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_44;
  wire       [6:0]    _zz_when_ArraySlice_l113_44;
  wire       [6:0]    _zz_when_ArraySlice_l113_44_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_44_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_44_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_44_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_44;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_44_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_44_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_44_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_44;
  wire       [6:0]    _zz_when_ArraySlice_l118_44_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_44_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_44_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_44_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_44_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_44_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_44_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_44_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_44_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_45;
  wire       [5:0]    _zz_when_ArraySlice_l165_45_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_45;
  wire       [4:0]    _zz_when_ArraySlice_l166_45_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_45_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_45_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_45_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_45;
  wire       [6:0]    _zz_when_ArraySlice_l113_45;
  wire       [6:0]    _zz_when_ArraySlice_l113_45_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_45_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_45_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_45_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_45;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_45_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_45_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_45_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_45;
  wire       [6:0]    _zz_when_ArraySlice_l118_45_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_45_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_45_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_45_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_45_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_45_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_45_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_45_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_45_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_46;
  wire       [5:0]    _zz_when_ArraySlice_l165_46_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_46;
  wire       [4:0]    _zz_when_ArraySlice_l166_46_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_46_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_46_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_46_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_46;
  wire       [6:0]    _zz_when_ArraySlice_l113_46;
  wire       [6:0]    _zz_when_ArraySlice_l113_46_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_46_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_46_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_46_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_46;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_46_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_46_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_46_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_46;
  wire       [6:0]    _zz_when_ArraySlice_l118_46_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_46_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_46_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_46_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_46_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_46_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_46_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_46_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_46_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_47;
  wire       [5:0]    _zz_when_ArraySlice_l165_47_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_47;
  wire       [3:0]    _zz_when_ArraySlice_l166_47_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_47_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_47_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_47_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_47;
  wire       [6:0]    _zz_when_ArraySlice_l113_47;
  wire       [6:0]    _zz_when_ArraySlice_l113_47_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_47_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_47_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_47_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_47;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_47_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_47_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_47_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_47;
  wire       [6:0]    _zz_when_ArraySlice_l118_47_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_47_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_47_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_47_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_47_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_47_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_47_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_47_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_47_8;
  wire                _zz_when_ArraySlice_l418_1_1;
  wire                _zz_when_ArraySlice_l418_1_2;
  wire                _zz_when_ArraySlice_l418_1_3;
  wire                _zz_when_ArraySlice_l418_1_4;
  wire                _zz_when_ArraySlice_l418_1_5;
  wire                _zz_when_ArraySlice_l418_1_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l421_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l421_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l421_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l421_1_5;
  wire       [0:0]    _zz_when_ArraySlice_l421_1_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_1_7;
  wire       [3:0]    _zz_when_ArraySlice_l421_1_8;
  wire       [5:0]    _zz_selectReadFifo_1_24;
  wire       [0:0]    _zz_selectReadFifo_1_25;
  wire       [12:0]   _zz_when_ArraySlice_l425_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l425_1_2;
  wire       [12:0]   _zz_when_ArraySlice_l425_1_3;
  wire       [0:0]    _zz_when_ArraySlice_l425_1_4;
  wire       [12:0]   _zz_when_ArraySlice_l436_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l436_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l436_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l436_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l436_1_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_5;
  wire       [6:0]    _zz_when_ArraySlice_l95_5;
  wire       [6:0]    _zz_when_ArraySlice_l95_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_5_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_5_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_1_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_1_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_1_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_5;
  wire       [6:0]    _zz_when_ArraySlice_l99_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_1_2;
  wire       [0:0]    _zz_when_ArraySlice_l437_1_3;
  wire       [6:0]    _zz_when_ArraySlice_l437_1_4;
  wire       [5:0]    _zz_selectReadFifo_1_26;
  wire       [5:0]    _zz_selectReadFifo_1_27;
  wire       [5:0]    _zz_selectReadFifo_1_28;
  wire       [0:0]    _zz_selectReadFifo_1_29;
  wire       [5:0]    _zz_when_ArraySlice_l165_48;
  wire       [5:0]    _zz_when_ArraySlice_l165_48_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_48_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_48;
  wire       [6:0]    _zz_when_ArraySlice_l166_48_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_48_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_48_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_48_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_48_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_48;
  wire       [6:0]    _zz_when_ArraySlice_l113_48;
  wire       [6:0]    _zz_when_ArraySlice_l113_48_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_48_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_48_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_48_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_48;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_48_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_48_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_48_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_48;
  wire       [6:0]    _zz_when_ArraySlice_l118_48_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_48_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_48_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_48_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_48_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_48_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_48_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_48_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_48_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_49;
  wire       [5:0]    _zz_when_ArraySlice_l165_49_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_49_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_49;
  wire       [5:0]    _zz_when_ArraySlice_l166_49_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_49_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_49_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_49_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_49;
  wire       [6:0]    _zz_when_ArraySlice_l113_49;
  wire       [6:0]    _zz_when_ArraySlice_l113_49_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_49_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_49_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_49_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_49;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_49_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_49_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_49_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_49;
  wire       [6:0]    _zz_when_ArraySlice_l118_49_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_49_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_49_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_49_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_49_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_49_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_49_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_49_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_49_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_49_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_50;
  wire       [5:0]    _zz_when_ArraySlice_l165_50_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_50_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_50;
  wire       [5:0]    _zz_when_ArraySlice_l166_50_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_50_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_50_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_50_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_50;
  wire       [6:0]    _zz_when_ArraySlice_l113_50;
  wire       [6:0]    _zz_when_ArraySlice_l113_50_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_50_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_50_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_50_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_50;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_50_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_50_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_50_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_50;
  wire       [6:0]    _zz_when_ArraySlice_l118_50_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_50_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_50_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_50_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_50_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_50_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_50_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_50_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_50_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_50_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_51;
  wire       [5:0]    _zz_when_ArraySlice_l165_51_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_51_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_51;
  wire       [5:0]    _zz_when_ArraySlice_l166_51_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_51_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_51_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_51_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_51;
  wire       [6:0]    _zz_when_ArraySlice_l113_51;
  wire       [6:0]    _zz_when_ArraySlice_l113_51_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_51_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_51_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_51_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_51;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_51_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_51_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_51_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_51;
  wire       [6:0]    _zz_when_ArraySlice_l118_51_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_51_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_51_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_51_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_51_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_51_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_51_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_51_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_51_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_51_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_52;
  wire       [5:0]    _zz_when_ArraySlice_l165_52_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_52;
  wire       [5:0]    _zz_when_ArraySlice_l166_52_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_52_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_52_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_52;
  wire       [6:0]    _zz_when_ArraySlice_l113_52;
  wire       [6:0]    _zz_when_ArraySlice_l113_52_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_52_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_52_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_52_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_52;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_52_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_52_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_52_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_52;
  wire       [6:0]    _zz_when_ArraySlice_l118_52_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_52_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_52_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_52_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_52_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_52_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_52_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_52_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_52_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_53;
  wire       [5:0]    _zz_when_ArraySlice_l165_53_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_53;
  wire       [4:0]    _zz_when_ArraySlice_l166_53_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_53_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_53_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_53_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_53;
  wire       [6:0]    _zz_when_ArraySlice_l113_53;
  wire       [6:0]    _zz_when_ArraySlice_l113_53_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_53_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_53_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_53_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_53;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_53_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_53_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_53_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_53;
  wire       [6:0]    _zz_when_ArraySlice_l118_53_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_53_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_53_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_53_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_53_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_53_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_53_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_53_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_53_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_54;
  wire       [5:0]    _zz_when_ArraySlice_l165_54_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_54;
  wire       [4:0]    _zz_when_ArraySlice_l166_54_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_54_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_54_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_54_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_54;
  wire       [6:0]    _zz_when_ArraySlice_l113_54;
  wire       [6:0]    _zz_when_ArraySlice_l113_54_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_54_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_54_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_54_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_54;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_54_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_54_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_54_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_54;
  wire       [6:0]    _zz_when_ArraySlice_l118_54_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_54_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_54_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_54_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_54_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_54_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_54_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_54_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_54_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_55;
  wire       [5:0]    _zz_when_ArraySlice_l165_55_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_55;
  wire       [3:0]    _zz_when_ArraySlice_l166_55_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_55_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_55_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_55_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_55;
  wire       [6:0]    _zz_when_ArraySlice_l113_55;
  wire       [6:0]    _zz_when_ArraySlice_l113_55_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_55_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_55_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_55_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_55;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_55_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_55_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_55_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_55;
  wire       [6:0]    _zz_when_ArraySlice_l118_55_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_55_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_55_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_55_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_55_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_55_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_55_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_55_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_55_8;
  wire                _zz_when_ArraySlice_l444_1_1;
  wire                _zz_when_ArraySlice_l444_1_2;
  wire                _zz_when_ArraySlice_l444_1_3;
  wire                _zz_when_ArraySlice_l444_1_4;
  wire                _zz_when_ArraySlice_l444_1_5;
  wire                _zz_when_ArraySlice_l444_1_6;
  wire       [5:0]    _zz_selectReadFifo_1_30;
  wire       [0:0]    _zz_selectReadFifo_1_31;
  wire       [12:0]   _zz_when_ArraySlice_l448_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l448_1_2;
  wire       [12:0]   _zz_when_ArraySlice_l448_1_3;
  wire       [0:0]    _zz_when_ArraySlice_l448_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l434_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l434_1_2;
  wire       [3:0]    _zz_when_ArraySlice_l434_1_3;
  wire       [12:0]   _zz_when_ArraySlice_l455_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l455_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l455_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l455_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l455_1_5;
  wire       [5:0]    _zz_when_ArraySlice_l373_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l373_2_2;
  wire       [4:0]    _zz_when_ArraySlice_l373_2_3;
  reg        [6:0]    _zz_when_ArraySlice_l374_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l374_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l374_2_3;
  wire       [4:0]    _zz_when_ArraySlice_l374_2_4;
  wire       [5:0]    _zz__zz_outputStreamArrayData_2_valid;
  wire       [4:0]    _zz__zz_outputStreamArrayData_2_valid_1;
  reg                 _zz_outputStreamArrayData_2_valid_2;
  reg        [31:0]   _zz_outputStreamArrayData_2_payload;
  wire       [6:0]    _zz_when_ArraySlice_l380_2_1;
  wire       [0:0]    _zz_when_ArraySlice_l380_2_2;
  reg        [6:0]    _zz_when_ArraySlice_l380_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l380_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l380_2_5;
  wire       [4:0]    _zz_when_ArraySlice_l380_2_6;
  wire       [12:0]   _zz_when_ArraySlice_l381_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l381_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l381_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l381_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l381_2_5;
  wire       [5:0]    _zz_selectReadFifo_2;
  wire       [5:0]    _zz_selectReadFifo_2_1;
  wire       [5:0]    _zz_selectReadFifo_2_2;
  wire       [0:0]    _zz_selectReadFifo_2_3;
  wire       [5:0]    _zz_selectReadFifo_2_4;
  wire       [0:0]    _zz_selectReadFifo_2_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_2_1;
  wire       [12:0]   _zz_when_ArraySlice_l384_2_2;
  wire       [12:0]   _zz_when_ArraySlice_l384_2_3;
  wire       [0:0]    _zz_when_ArraySlice_l384_2_4;
  reg        [6:0]    _zz_when_ArraySlice_l389_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l389_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l389_2_3;
  wire       [4:0]    _zz_when_ArraySlice_l389_2_4;
  wire       [6:0]    _zz_when_ArraySlice_l389_2_5;
  wire       [0:0]    _zz_when_ArraySlice_l389_2_6;
  wire       [12:0]   _zz_when_ArraySlice_l390_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l390_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l390_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l390_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l390_2_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_6;
  wire       [6:0]    _zz_when_ArraySlice_l95_6;
  wire       [6:0]    _zz_when_ArraySlice_l95_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_6_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_6_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_2_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_2_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_2_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_6;
  wire       [6:0]    _zz_when_ArraySlice_l99_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_2_2;
  wire       [0:0]    _zz_when_ArraySlice_l392_2_3;
  wire       [6:0]    _zz_when_ArraySlice_l392_2_4;
  wire       [5:0]    _zz_selectReadFifo_2_6;
  wire       [5:0]    _zz_selectReadFifo_2_7;
  wire       [5:0]    _zz_selectReadFifo_2_8;
  wire       [0:0]    _zz_selectReadFifo_2_9;
  wire       [5:0]    _zz_selectReadFifo_2_10;
  wire       [5:0]    _zz_selectReadFifo_2_11;
  wire       [5:0]    _zz_selectReadFifo_2_12;
  wire       [0:0]    _zz_selectReadFifo_2_13;
  wire       [5:0]    _zz_when_ArraySlice_l165_56;
  wire       [5:0]    _zz_when_ArraySlice_l165_56_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_56_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_56;
  wire       [6:0]    _zz_when_ArraySlice_l166_56_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_56_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_56_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_56_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_56_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_56;
  wire       [6:0]    _zz_when_ArraySlice_l113_56;
  wire       [6:0]    _zz_when_ArraySlice_l113_56_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_56_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_56_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_56_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_56;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_56_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_56_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_56_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_56;
  wire       [6:0]    _zz_when_ArraySlice_l118_56_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_56_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_56_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_56_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_56_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_56_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_56_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_56_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_56_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_57;
  wire       [5:0]    _zz_when_ArraySlice_l165_57_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_57_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_57;
  wire       [5:0]    _zz_when_ArraySlice_l166_57_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_57_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_57_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_57_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_57;
  wire       [6:0]    _zz_when_ArraySlice_l113_57;
  wire       [6:0]    _zz_when_ArraySlice_l113_57_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_57_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_57_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_57_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_57;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_57_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_57_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_57_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_57;
  wire       [6:0]    _zz_when_ArraySlice_l118_57_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_57_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_57_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_57_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_57_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_57_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_57_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_57_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_57_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_57_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_58;
  wire       [5:0]    _zz_when_ArraySlice_l165_58_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_58_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_58;
  wire       [5:0]    _zz_when_ArraySlice_l166_58_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_58_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_58_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_58_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_58;
  wire       [6:0]    _zz_when_ArraySlice_l113_58;
  wire       [6:0]    _zz_when_ArraySlice_l113_58_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_58_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_58_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_58_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_58;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_58_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_58_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_58_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_58;
  wire       [6:0]    _zz_when_ArraySlice_l118_58_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_58_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_58_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_58_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_58_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_58_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_58_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_58_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_58_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_58_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_59;
  wire       [5:0]    _zz_when_ArraySlice_l165_59_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_59_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_59;
  wire       [5:0]    _zz_when_ArraySlice_l166_59_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_59_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_59_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_59_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_59;
  wire       [6:0]    _zz_when_ArraySlice_l113_59;
  wire       [6:0]    _zz_when_ArraySlice_l113_59_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_59_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_59_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_59_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_59;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_59_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_59_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_59_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_59;
  wire       [6:0]    _zz_when_ArraySlice_l118_59_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_59_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_59_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_59_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_59_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_59_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_59_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_59_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_59_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_59_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_60;
  wire       [5:0]    _zz_when_ArraySlice_l165_60_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_60;
  wire       [5:0]    _zz_when_ArraySlice_l166_60_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_60_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_60_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_60;
  wire       [6:0]    _zz_when_ArraySlice_l113_60;
  wire       [6:0]    _zz_when_ArraySlice_l113_60_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_60_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_60_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_60_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_60;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_60_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_60_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_60_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_60;
  wire       [6:0]    _zz_when_ArraySlice_l118_60_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_60_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_60_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_60_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_60_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_60_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_60_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_60_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_60_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_61;
  wire       [5:0]    _zz_when_ArraySlice_l165_61_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_61;
  wire       [4:0]    _zz_when_ArraySlice_l166_61_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_61_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_61_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_61_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_61;
  wire       [6:0]    _zz_when_ArraySlice_l113_61;
  wire       [6:0]    _zz_when_ArraySlice_l113_61_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_61_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_61_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_61_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_61;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_61_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_61_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_61_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_61;
  wire       [6:0]    _zz_when_ArraySlice_l118_61_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_61_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_61_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_61_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_61_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_61_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_61_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_61_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_61_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_62;
  wire       [5:0]    _zz_when_ArraySlice_l165_62_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_62;
  wire       [4:0]    _zz_when_ArraySlice_l166_62_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_62_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_62_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_62_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_62;
  wire       [6:0]    _zz_when_ArraySlice_l113_62;
  wire       [6:0]    _zz_when_ArraySlice_l113_62_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_62_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_62_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_62_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_62;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_62_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_62_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_62_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_62;
  wire       [6:0]    _zz_when_ArraySlice_l118_62_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_62_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_62_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_62_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_62_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_62_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_62_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_62_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_62_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_63;
  wire       [5:0]    _zz_when_ArraySlice_l165_63_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_63;
  wire       [3:0]    _zz_when_ArraySlice_l166_63_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_63_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_63_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_63_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_63;
  wire       [6:0]    _zz_when_ArraySlice_l113_63;
  wire       [6:0]    _zz_when_ArraySlice_l113_63_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_63_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_63_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_63_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_63;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_63_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_63_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_63_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_63;
  wire       [6:0]    _zz_when_ArraySlice_l118_63_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_63_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_63_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_63_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_63_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_63_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_63_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_63_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_63_8;
  wire                _zz_when_ArraySlice_l398_2_1;
  wire                _zz_when_ArraySlice_l398_2_2;
  wire                _zz_when_ArraySlice_l398_2_3;
  wire                _zz_when_ArraySlice_l398_2_4;
  wire                _zz_when_ArraySlice_l398_2_5;
  wire                _zz_when_ArraySlice_l398_2_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l401_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l401_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l401_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l401_2_5;
  wire       [0:0]    _zz_when_ArraySlice_l401_2_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_2_7;
  wire       [4:0]    _zz_when_ArraySlice_l401_2_8;
  wire       [5:0]    _zz_selectReadFifo_2_14;
  wire       [0:0]    _zz_selectReadFifo_2_15;
  wire       [12:0]   _zz_when_ArraySlice_l405_2_1;
  wire       [12:0]   _zz_when_ArraySlice_l405_2_2;
  wire       [12:0]   _zz_when_ArraySlice_l405_2_3;
  wire       [0:0]    _zz_when_ArraySlice_l405_2_4;
  reg        [6:0]    _zz_when_ArraySlice_l409_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l409_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l409_2_3;
  wire       [4:0]    _zz_when_ArraySlice_l409_2_4;
  wire       [12:0]   _zz_when_ArraySlice_l410_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l410_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l410_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l410_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l410_2_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_7;
  wire       [6:0]    _zz_when_ArraySlice_l95_7;
  wire       [6:0]    _zz_when_ArraySlice_l95_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_7_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_7_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_2_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_2_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_2_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_7;
  wire       [6:0]    _zz_when_ArraySlice_l99_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_2_2;
  wire       [0:0]    _zz_when_ArraySlice_l412_2_3;
  wire       [6:0]    _zz_when_ArraySlice_l412_2_4;
  wire       [5:0]    _zz_selectReadFifo_2_16;
  wire       [5:0]    _zz_selectReadFifo_2_17;
  wire       [5:0]    _zz_selectReadFifo_2_18;
  wire       [0:0]    _zz_selectReadFifo_2_19;
  wire       [5:0]    _zz_selectReadFifo_2_20;
  wire       [5:0]    _zz_selectReadFifo_2_21;
  wire       [5:0]    _zz_selectReadFifo_2_22;
  wire       [0:0]    _zz_selectReadFifo_2_23;
  wire       [5:0]    _zz_when_ArraySlice_l165_64;
  wire       [5:0]    _zz_when_ArraySlice_l165_64_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_64_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_64;
  wire       [6:0]    _zz_when_ArraySlice_l166_64_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_64_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_64_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_64_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_64_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_64;
  wire       [6:0]    _zz_when_ArraySlice_l113_64;
  wire       [6:0]    _zz_when_ArraySlice_l113_64_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_64_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_64_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_64_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_64;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_64_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_64_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_64_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_64;
  wire       [6:0]    _zz_when_ArraySlice_l118_64_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_64_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_64_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_64_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_64_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_64_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_64_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_64_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_64_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_65;
  wire       [5:0]    _zz_when_ArraySlice_l165_65_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_65_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_65;
  wire       [5:0]    _zz_when_ArraySlice_l166_65_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_65_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_65_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_65_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_65;
  wire       [6:0]    _zz_when_ArraySlice_l113_65;
  wire       [6:0]    _zz_when_ArraySlice_l113_65_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_65_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_65_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_65_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_65;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_65_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_65_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_65_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_65;
  wire       [6:0]    _zz_when_ArraySlice_l118_65_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_65_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_65_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_65_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_65_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_65_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_65_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_65_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_65_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_65_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_66;
  wire       [5:0]    _zz_when_ArraySlice_l165_66_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_66_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_66;
  wire       [5:0]    _zz_when_ArraySlice_l166_66_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_66_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_66_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_66_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_66;
  wire       [6:0]    _zz_when_ArraySlice_l113_66;
  wire       [6:0]    _zz_when_ArraySlice_l113_66_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_66_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_66_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_66_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_66;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_66_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_66_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_66_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_66;
  wire       [6:0]    _zz_when_ArraySlice_l118_66_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_66_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_66_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_66_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_66_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_66_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_66_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_66_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_66_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_66_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_67;
  wire       [5:0]    _zz_when_ArraySlice_l165_67_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_67_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_67;
  wire       [5:0]    _zz_when_ArraySlice_l166_67_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_67_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_67_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_67_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_67;
  wire       [6:0]    _zz_when_ArraySlice_l113_67;
  wire       [6:0]    _zz_when_ArraySlice_l113_67_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_67_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_67_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_67_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_67;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_67_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_67_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_67_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_67;
  wire       [6:0]    _zz_when_ArraySlice_l118_67_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_67_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_67_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_67_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_67_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_67_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_67_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_67_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_67_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_67_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_68;
  wire       [5:0]    _zz_when_ArraySlice_l165_68_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_68;
  wire       [5:0]    _zz_when_ArraySlice_l166_68_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_68_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_68_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_68;
  wire       [6:0]    _zz_when_ArraySlice_l113_68;
  wire       [6:0]    _zz_when_ArraySlice_l113_68_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_68_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_68_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_68_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_68;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_68_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_68_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_68_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_68;
  wire       [6:0]    _zz_when_ArraySlice_l118_68_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_68_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_68_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_68_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_68_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_68_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_68_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_68_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_68_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_69;
  wire       [5:0]    _zz_when_ArraySlice_l165_69_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_69;
  wire       [4:0]    _zz_when_ArraySlice_l166_69_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_69_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_69_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_69_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_69;
  wire       [6:0]    _zz_when_ArraySlice_l113_69;
  wire       [6:0]    _zz_when_ArraySlice_l113_69_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_69_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_69_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_69_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_69;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_69_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_69_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_69_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_69;
  wire       [6:0]    _zz_when_ArraySlice_l118_69_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_69_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_69_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_69_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_69_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_69_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_69_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_69_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_69_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_70;
  wire       [5:0]    _zz_when_ArraySlice_l165_70_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_70;
  wire       [4:0]    _zz_when_ArraySlice_l166_70_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_70_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_70_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_70_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_70;
  wire       [6:0]    _zz_when_ArraySlice_l113_70;
  wire       [6:0]    _zz_when_ArraySlice_l113_70_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_70_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_70_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_70_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_70;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_70_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_70_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_70_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_70;
  wire       [6:0]    _zz_when_ArraySlice_l118_70_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_70_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_70_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_70_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_70_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_70_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_70_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_70_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_70_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_71;
  wire       [5:0]    _zz_when_ArraySlice_l165_71_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_71;
  wire       [3:0]    _zz_when_ArraySlice_l166_71_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_71_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_71_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_71_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_71;
  wire       [6:0]    _zz_when_ArraySlice_l113_71;
  wire       [6:0]    _zz_when_ArraySlice_l113_71_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_71_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_71_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_71_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_71;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_71_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_71_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_71_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_71;
  wire       [6:0]    _zz_when_ArraySlice_l118_71_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_71_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_71_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_71_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_71_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_71_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_71_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_71_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_71_8;
  wire                _zz_when_ArraySlice_l418_2_1;
  wire                _zz_when_ArraySlice_l418_2_2;
  wire                _zz_when_ArraySlice_l418_2_3;
  wire                _zz_when_ArraySlice_l418_2_4;
  wire                _zz_when_ArraySlice_l418_2_5;
  wire                _zz_when_ArraySlice_l418_2_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l421_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l421_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l421_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l421_2_5;
  wire       [0:0]    _zz_when_ArraySlice_l421_2_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_2_7;
  wire       [4:0]    _zz_when_ArraySlice_l421_2_8;
  wire       [5:0]    _zz_selectReadFifo_2_24;
  wire       [0:0]    _zz_selectReadFifo_2_25;
  wire       [12:0]   _zz_when_ArraySlice_l425_2_1;
  wire       [12:0]   _zz_when_ArraySlice_l425_2_2;
  wire       [12:0]   _zz_when_ArraySlice_l425_2_3;
  wire       [0:0]    _zz_when_ArraySlice_l425_2_4;
  wire       [12:0]   _zz_when_ArraySlice_l436_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l436_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l436_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l436_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l436_2_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_8;
  wire       [6:0]    _zz_when_ArraySlice_l95_8;
  wire       [6:0]    _zz_when_ArraySlice_l95_8_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_8_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_8_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_8_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_2_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_2_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_2_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_8;
  wire       [6:0]    _zz_when_ArraySlice_l99_8_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_2_2;
  wire       [0:0]    _zz_when_ArraySlice_l437_2_3;
  wire       [6:0]    _zz_when_ArraySlice_l437_2_4;
  wire       [5:0]    _zz_selectReadFifo_2_26;
  wire       [5:0]    _zz_selectReadFifo_2_27;
  wire       [5:0]    _zz_selectReadFifo_2_28;
  wire       [0:0]    _zz_selectReadFifo_2_29;
  wire       [5:0]    _zz_when_ArraySlice_l165_72;
  wire       [5:0]    _zz_when_ArraySlice_l165_72_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_72_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_72;
  wire       [6:0]    _zz_when_ArraySlice_l166_72_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_72_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_72_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_72_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_72_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_72;
  wire       [6:0]    _zz_when_ArraySlice_l113_72;
  wire       [6:0]    _zz_when_ArraySlice_l113_72_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_72_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_72_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_72_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_72;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_72_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_72_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_72_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_72;
  wire       [6:0]    _zz_when_ArraySlice_l118_72_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_72_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_72_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_72_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_72_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_72_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_72_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_72_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_72_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_73;
  wire       [5:0]    _zz_when_ArraySlice_l165_73_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_73_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_73;
  wire       [5:0]    _zz_when_ArraySlice_l166_73_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_73_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_73_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_73_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_73;
  wire       [6:0]    _zz_when_ArraySlice_l113_73;
  wire       [6:0]    _zz_when_ArraySlice_l113_73_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_73_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_73_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_73_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_73;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_73_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_73_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_73_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_73;
  wire       [6:0]    _zz_when_ArraySlice_l118_73_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_73_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_73_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_73_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_73_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_73_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_73_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_73_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_73_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_73_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_74;
  wire       [5:0]    _zz_when_ArraySlice_l165_74_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_74_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_74;
  wire       [5:0]    _zz_when_ArraySlice_l166_74_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_74_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_74_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_74_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_74;
  wire       [6:0]    _zz_when_ArraySlice_l113_74;
  wire       [6:0]    _zz_when_ArraySlice_l113_74_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_74_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_74_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_74_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_74;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_74_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_74_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_74_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_74;
  wire       [6:0]    _zz_when_ArraySlice_l118_74_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_74_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_74_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_74_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_74_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_74_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_74_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_74_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_74_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_74_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_75;
  wire       [5:0]    _zz_when_ArraySlice_l165_75_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_75_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_75;
  wire       [5:0]    _zz_when_ArraySlice_l166_75_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_75_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_75_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_75_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_75;
  wire       [6:0]    _zz_when_ArraySlice_l113_75;
  wire       [6:0]    _zz_when_ArraySlice_l113_75_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_75_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_75_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_75_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_75;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_75_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_75_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_75_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_75;
  wire       [6:0]    _zz_when_ArraySlice_l118_75_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_75_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_75_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_75_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_75_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_75_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_75_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_75_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_75_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_75_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_76;
  wire       [5:0]    _zz_when_ArraySlice_l165_76_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_76;
  wire       [5:0]    _zz_when_ArraySlice_l166_76_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_76_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_76_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_76;
  wire       [6:0]    _zz_when_ArraySlice_l113_76;
  wire       [6:0]    _zz_when_ArraySlice_l113_76_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_76_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_76_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_76_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_76;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_76_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_76_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_76_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_76;
  wire       [6:0]    _zz_when_ArraySlice_l118_76_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_76_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_76_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_76_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_76_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_76_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_76_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_76_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_76_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_77;
  wire       [5:0]    _zz_when_ArraySlice_l165_77_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_77;
  wire       [4:0]    _zz_when_ArraySlice_l166_77_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_77_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_77_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_77_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_77;
  wire       [6:0]    _zz_when_ArraySlice_l113_77;
  wire       [6:0]    _zz_when_ArraySlice_l113_77_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_77_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_77_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_77_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_77;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_77_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_77_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_77_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_77;
  wire       [6:0]    _zz_when_ArraySlice_l118_77_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_77_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_77_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_77_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_77_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_77_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_77_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_77_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_77_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_78;
  wire       [5:0]    _zz_when_ArraySlice_l165_78_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_78;
  wire       [4:0]    _zz_when_ArraySlice_l166_78_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_78_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_78_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_78_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_78;
  wire       [6:0]    _zz_when_ArraySlice_l113_78;
  wire       [6:0]    _zz_when_ArraySlice_l113_78_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_78_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_78_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_78_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_78;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_78_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_78_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_78_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_78;
  wire       [6:0]    _zz_when_ArraySlice_l118_78_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_78_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_78_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_78_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_78_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_78_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_78_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_78_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_78_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_79;
  wire       [5:0]    _zz_when_ArraySlice_l165_79_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_79;
  wire       [3:0]    _zz_when_ArraySlice_l166_79_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_79_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_79_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_79_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_79;
  wire       [6:0]    _zz_when_ArraySlice_l113_79;
  wire       [6:0]    _zz_when_ArraySlice_l113_79_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_79_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_79_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_79_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_79;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_79_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_79_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_79_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_79;
  wire       [6:0]    _zz_when_ArraySlice_l118_79_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_79_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_79_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_79_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_79_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_79_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_79_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_79_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_79_8;
  wire                _zz_when_ArraySlice_l444_2_1;
  wire                _zz_when_ArraySlice_l444_2_2;
  wire                _zz_when_ArraySlice_l444_2_3;
  wire                _zz_when_ArraySlice_l444_2_4;
  wire                _zz_when_ArraySlice_l444_2_5;
  wire                _zz_when_ArraySlice_l444_2_6;
  wire       [5:0]    _zz_selectReadFifo_2_30;
  wire       [0:0]    _zz_selectReadFifo_2_31;
  wire       [12:0]   _zz_when_ArraySlice_l448_2_1;
  wire       [12:0]   _zz_when_ArraySlice_l448_2_2;
  wire       [12:0]   _zz_when_ArraySlice_l448_2_3;
  wire       [0:0]    _zz_when_ArraySlice_l448_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l434_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l434_2_2;
  wire       [4:0]    _zz_when_ArraySlice_l434_2_3;
  wire       [12:0]   _zz_when_ArraySlice_l455_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l455_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l455_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l455_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l455_2_5;
  wire       [5:0]    _zz_when_ArraySlice_l373_3;
  wire       [5:0]    _zz_when_ArraySlice_l373_3_1;
  wire       [4:0]    _zz_when_ArraySlice_l373_3_2;
  reg        [6:0]    _zz_when_ArraySlice_l374_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l374_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l374_3_3;
  wire       [4:0]    _zz_when_ArraySlice_l374_3_4;
  wire       [5:0]    _zz__zz_outputStreamArrayData_3_valid;
  wire       [4:0]    _zz__zz_outputStreamArrayData_3_valid_1;
  reg                 _zz_outputStreamArrayData_3_valid_2;
  reg        [31:0]   _zz_outputStreamArrayData_3_payload;
  wire       [6:0]    _zz_when_ArraySlice_l380_3_1;
  wire       [0:0]    _zz_when_ArraySlice_l380_3_2;
  reg        [6:0]    _zz_when_ArraySlice_l380_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l380_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l380_3_5;
  wire       [4:0]    _zz_when_ArraySlice_l380_3_6;
  wire       [12:0]   _zz_when_ArraySlice_l381_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l381_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l381_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l381_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l381_3_5;
  wire       [5:0]    _zz_selectReadFifo_3;
  wire       [5:0]    _zz_selectReadFifo_3_1;
  wire       [5:0]    _zz_selectReadFifo_3_2;
  wire       [0:0]    _zz_selectReadFifo_3_3;
  wire       [5:0]    _zz_selectReadFifo_3_4;
  wire       [0:0]    _zz_selectReadFifo_3_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_3_1;
  wire       [12:0]   _zz_when_ArraySlice_l384_3_2;
  wire       [12:0]   _zz_when_ArraySlice_l384_3_3;
  wire       [0:0]    _zz_when_ArraySlice_l384_3_4;
  reg        [6:0]    _zz_when_ArraySlice_l389_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l389_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l389_3_3;
  wire       [4:0]    _zz_when_ArraySlice_l389_3_4;
  wire       [6:0]    _zz_when_ArraySlice_l389_3_5;
  wire       [0:0]    _zz_when_ArraySlice_l389_3_6;
  wire       [12:0]   _zz_when_ArraySlice_l390_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l390_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l390_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l390_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l390_3_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_9;
  wire       [6:0]    _zz_when_ArraySlice_l95_9;
  wire       [6:0]    _zz_when_ArraySlice_l95_9_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_9_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_9_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_9_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_3_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_3_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_3_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_9;
  wire       [6:0]    _zz_when_ArraySlice_l99_9_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_3_2;
  wire       [0:0]    _zz_when_ArraySlice_l392_3_3;
  wire       [6:0]    _zz_when_ArraySlice_l392_3_4;
  wire       [5:0]    _zz_selectReadFifo_3_6;
  wire       [5:0]    _zz_selectReadFifo_3_7;
  wire       [5:0]    _zz_selectReadFifo_3_8;
  wire       [0:0]    _zz_selectReadFifo_3_9;
  wire       [5:0]    _zz_selectReadFifo_3_10;
  wire       [5:0]    _zz_selectReadFifo_3_11;
  wire       [5:0]    _zz_selectReadFifo_3_12;
  wire       [0:0]    _zz_selectReadFifo_3_13;
  wire       [5:0]    _zz_when_ArraySlice_l165_80;
  wire       [5:0]    _zz_when_ArraySlice_l165_80_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_80_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_80;
  wire       [6:0]    _zz_when_ArraySlice_l166_80_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_80_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_80_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_80_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_80_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_80;
  wire       [6:0]    _zz_when_ArraySlice_l113_80;
  wire       [6:0]    _zz_when_ArraySlice_l113_80_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_80_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_80_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_80_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_80;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_80_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_80_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_80_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_80;
  wire       [6:0]    _zz_when_ArraySlice_l118_80_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_80_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_80_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_80_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_80_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_80_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_80_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_80_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_80_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_81;
  wire       [5:0]    _zz_when_ArraySlice_l165_81_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_81_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_81;
  wire       [5:0]    _zz_when_ArraySlice_l166_81_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_81_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_81_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_81_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_81;
  wire       [6:0]    _zz_when_ArraySlice_l113_81;
  wire       [6:0]    _zz_when_ArraySlice_l113_81_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_81_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_81_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_81_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_81;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_81_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_81_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_81_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_81;
  wire       [6:0]    _zz_when_ArraySlice_l118_81_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_81_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_81_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_81_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_81_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_81_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_81_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_81_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_81_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_81_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_82;
  wire       [5:0]    _zz_when_ArraySlice_l165_82_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_82_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_82;
  wire       [5:0]    _zz_when_ArraySlice_l166_82_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_82_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_82_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_82_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_82;
  wire       [6:0]    _zz_when_ArraySlice_l113_82;
  wire       [6:0]    _zz_when_ArraySlice_l113_82_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_82_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_82_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_82_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_82;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_82_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_82_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_82_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_82;
  wire       [6:0]    _zz_when_ArraySlice_l118_82_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_82_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_82_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_82_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_82_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_82_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_82_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_82_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_82_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_82_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_83;
  wire       [5:0]    _zz_when_ArraySlice_l165_83_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_83_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_83;
  wire       [5:0]    _zz_when_ArraySlice_l166_83_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_83_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_83_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_83_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_83;
  wire       [6:0]    _zz_when_ArraySlice_l113_83;
  wire       [6:0]    _zz_when_ArraySlice_l113_83_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_83_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_83_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_83_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_83;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_83_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_83_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_83_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_83;
  wire       [6:0]    _zz_when_ArraySlice_l118_83_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_83_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_83_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_83_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_83_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_83_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_83_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_83_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_83_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_83_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_84;
  wire       [5:0]    _zz_when_ArraySlice_l165_84_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_84;
  wire       [5:0]    _zz_when_ArraySlice_l166_84_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_84_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_84_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_84;
  wire       [6:0]    _zz_when_ArraySlice_l113_84;
  wire       [6:0]    _zz_when_ArraySlice_l113_84_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_84_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_84_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_84_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_84;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_84_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_84_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_84_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_84;
  wire       [6:0]    _zz_when_ArraySlice_l118_84_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_84_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_84_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_84_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_84_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_84_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_84_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_84_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_84_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_85;
  wire       [5:0]    _zz_when_ArraySlice_l165_85_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_85;
  wire       [4:0]    _zz_when_ArraySlice_l166_85_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_85_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_85_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_85_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_85;
  wire       [6:0]    _zz_when_ArraySlice_l113_85;
  wire       [6:0]    _zz_when_ArraySlice_l113_85_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_85_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_85_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_85_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_85;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_85_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_85_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_85_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_85;
  wire       [6:0]    _zz_when_ArraySlice_l118_85_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_85_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_85_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_85_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_85_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_85_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_85_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_85_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_85_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_86;
  wire       [5:0]    _zz_when_ArraySlice_l165_86_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_86;
  wire       [4:0]    _zz_when_ArraySlice_l166_86_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_86_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_86_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_86_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_86;
  wire       [6:0]    _zz_when_ArraySlice_l113_86;
  wire       [6:0]    _zz_when_ArraySlice_l113_86_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_86_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_86_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_86_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_86;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_86_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_86_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_86_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_86;
  wire       [6:0]    _zz_when_ArraySlice_l118_86_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_86_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_86_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_86_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_86_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_86_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_86_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_86_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_86_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_87;
  wire       [5:0]    _zz_when_ArraySlice_l165_87_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_87;
  wire       [3:0]    _zz_when_ArraySlice_l166_87_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_87_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_87_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_87_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_87;
  wire       [6:0]    _zz_when_ArraySlice_l113_87;
  wire       [6:0]    _zz_when_ArraySlice_l113_87_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_87_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_87_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_87_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_87;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_87_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_87_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_87_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_87;
  wire       [6:0]    _zz_when_ArraySlice_l118_87_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_87_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_87_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_87_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_87_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_87_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_87_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_87_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_87_8;
  wire                _zz_when_ArraySlice_l398_3_1;
  wire                _zz_when_ArraySlice_l398_3_2;
  wire                _zz_when_ArraySlice_l398_3_3;
  wire                _zz_when_ArraySlice_l398_3_4;
  wire                _zz_when_ArraySlice_l398_3_5;
  wire                _zz_when_ArraySlice_l398_3_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l401_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l401_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l401_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l401_3_5;
  wire       [0:0]    _zz_when_ArraySlice_l401_3_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_3_7;
  wire       [4:0]    _zz_when_ArraySlice_l401_3_8;
  wire       [5:0]    _zz_selectReadFifo_3_14;
  wire       [0:0]    _zz_selectReadFifo_3_15;
  wire       [12:0]   _zz_when_ArraySlice_l405_3_1;
  wire       [12:0]   _zz_when_ArraySlice_l405_3_2;
  wire       [12:0]   _zz_when_ArraySlice_l405_3_3;
  wire       [0:0]    _zz_when_ArraySlice_l405_3_4;
  reg        [6:0]    _zz_when_ArraySlice_l409_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l409_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l409_3_3;
  wire       [4:0]    _zz_when_ArraySlice_l409_3_4;
  wire       [12:0]   _zz_when_ArraySlice_l410_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l410_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l410_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l410_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l410_3_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_10;
  wire       [6:0]    _zz_when_ArraySlice_l95_10;
  wire       [6:0]    _zz_when_ArraySlice_l95_10_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_10_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_10_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_10_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_3_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_3_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_3_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_10;
  wire       [6:0]    _zz_when_ArraySlice_l99_10_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_3_2;
  wire       [0:0]    _zz_when_ArraySlice_l412_3_3;
  wire       [6:0]    _zz_when_ArraySlice_l412_3_4;
  wire       [5:0]    _zz_selectReadFifo_3_16;
  wire       [5:0]    _zz_selectReadFifo_3_17;
  wire       [5:0]    _zz_selectReadFifo_3_18;
  wire       [0:0]    _zz_selectReadFifo_3_19;
  wire       [5:0]    _zz_selectReadFifo_3_20;
  wire       [5:0]    _zz_selectReadFifo_3_21;
  wire       [5:0]    _zz_selectReadFifo_3_22;
  wire       [0:0]    _zz_selectReadFifo_3_23;
  wire       [5:0]    _zz_when_ArraySlice_l165_88;
  wire       [5:0]    _zz_when_ArraySlice_l165_88_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_88_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_88;
  wire       [6:0]    _zz_when_ArraySlice_l166_88_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_88_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_88_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_88_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_88_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_88;
  wire       [6:0]    _zz_when_ArraySlice_l113_88;
  wire       [6:0]    _zz_when_ArraySlice_l113_88_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_88_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_88_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_88_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_88;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_88_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_88_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_88_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_88;
  wire       [6:0]    _zz_when_ArraySlice_l118_88_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_88_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_88_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_88_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_88_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_88_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_88_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_88_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_88_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_89;
  wire       [5:0]    _zz_when_ArraySlice_l165_89_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_89_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_89;
  wire       [5:0]    _zz_when_ArraySlice_l166_89_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_89_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_89_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_89_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_89;
  wire       [6:0]    _zz_when_ArraySlice_l113_89;
  wire       [6:0]    _zz_when_ArraySlice_l113_89_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_89_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_89_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_89_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_89;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_89_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_89_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_89_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_89;
  wire       [6:0]    _zz_when_ArraySlice_l118_89_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_89_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_89_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_89_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_89_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_89_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_89_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_89_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_89_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_89_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_90;
  wire       [5:0]    _zz_when_ArraySlice_l165_90_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_90_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_90;
  wire       [5:0]    _zz_when_ArraySlice_l166_90_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_90_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_90_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_90_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_90;
  wire       [6:0]    _zz_when_ArraySlice_l113_90;
  wire       [6:0]    _zz_when_ArraySlice_l113_90_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_90_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_90_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_90_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_90;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_90_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_90_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_90_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_90;
  wire       [6:0]    _zz_when_ArraySlice_l118_90_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_90_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_90_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_90_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_90_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_90_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_90_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_90_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_90_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_90_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_91;
  wire       [5:0]    _zz_when_ArraySlice_l165_91_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_91_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_91;
  wire       [5:0]    _zz_when_ArraySlice_l166_91_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_91_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_91_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_91_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_91;
  wire       [6:0]    _zz_when_ArraySlice_l113_91;
  wire       [6:0]    _zz_when_ArraySlice_l113_91_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_91_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_91_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_91_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_91;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_91_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_91_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_91_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_91;
  wire       [6:0]    _zz_when_ArraySlice_l118_91_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_91_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_91_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_91_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_91_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_91_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_91_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_91_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_91_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_91_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_92;
  wire       [5:0]    _zz_when_ArraySlice_l165_92_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_92;
  wire       [5:0]    _zz_when_ArraySlice_l166_92_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_92_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_92_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_92;
  wire       [6:0]    _zz_when_ArraySlice_l113_92;
  wire       [6:0]    _zz_when_ArraySlice_l113_92_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_92_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_92_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_92_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_92;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_92_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_92_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_92_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_92;
  wire       [6:0]    _zz_when_ArraySlice_l118_92_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_92_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_92_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_92_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_92_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_92_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_92_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_92_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_92_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_93;
  wire       [5:0]    _zz_when_ArraySlice_l165_93_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_93;
  wire       [4:0]    _zz_when_ArraySlice_l166_93_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_93_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_93_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_93_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_93;
  wire       [6:0]    _zz_when_ArraySlice_l113_93;
  wire       [6:0]    _zz_when_ArraySlice_l113_93_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_93_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_93_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_93_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_93;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_93_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_93_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_93_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_93;
  wire       [6:0]    _zz_when_ArraySlice_l118_93_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_93_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_93_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_93_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_93_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_93_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_93_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_93_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_93_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_94;
  wire       [5:0]    _zz_when_ArraySlice_l165_94_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_94;
  wire       [4:0]    _zz_when_ArraySlice_l166_94_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_94_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_94_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_94_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_94;
  wire       [6:0]    _zz_when_ArraySlice_l113_94;
  wire       [6:0]    _zz_when_ArraySlice_l113_94_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_94_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_94_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_94_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_94;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_94_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_94_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_94_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_94;
  wire       [6:0]    _zz_when_ArraySlice_l118_94_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_94_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_94_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_94_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_94_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_94_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_94_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_94_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_94_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_95;
  wire       [5:0]    _zz_when_ArraySlice_l165_95_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_95;
  wire       [3:0]    _zz_when_ArraySlice_l166_95_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_95_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_95_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_95_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_95;
  wire       [6:0]    _zz_when_ArraySlice_l113_95;
  wire       [6:0]    _zz_when_ArraySlice_l113_95_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_95_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_95_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_95_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_95;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_95_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_95_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_95_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_95;
  wire       [6:0]    _zz_when_ArraySlice_l118_95_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_95_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_95_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_95_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_95_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_95_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_95_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_95_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_95_8;
  wire                _zz_when_ArraySlice_l418_3_1;
  wire                _zz_when_ArraySlice_l418_3_2;
  wire                _zz_when_ArraySlice_l418_3_3;
  wire                _zz_when_ArraySlice_l418_3_4;
  wire                _zz_when_ArraySlice_l418_3_5;
  wire                _zz_when_ArraySlice_l418_3_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l421_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l421_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l421_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l421_3_5;
  wire       [0:0]    _zz_when_ArraySlice_l421_3_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_3_7;
  wire       [4:0]    _zz_when_ArraySlice_l421_3_8;
  wire       [5:0]    _zz_selectReadFifo_3_24;
  wire       [0:0]    _zz_selectReadFifo_3_25;
  wire       [12:0]   _zz_when_ArraySlice_l425_3_1;
  wire       [12:0]   _zz_when_ArraySlice_l425_3_2;
  wire       [12:0]   _zz_when_ArraySlice_l425_3_3;
  wire       [0:0]    _zz_when_ArraySlice_l425_3_4;
  wire       [12:0]   _zz_when_ArraySlice_l436_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l436_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l436_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l436_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l436_3_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_11;
  wire       [6:0]    _zz_when_ArraySlice_l95_11;
  wire       [6:0]    _zz_when_ArraySlice_l95_11_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_11_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_11_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_11_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_3_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_3_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_3_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_11;
  wire       [6:0]    _zz_when_ArraySlice_l99_11_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_3_2;
  wire       [0:0]    _zz_when_ArraySlice_l437_3_3;
  wire       [6:0]    _zz_when_ArraySlice_l437_3_4;
  wire       [5:0]    _zz_selectReadFifo_3_26;
  wire       [5:0]    _zz_selectReadFifo_3_27;
  wire       [5:0]    _zz_selectReadFifo_3_28;
  wire       [0:0]    _zz_selectReadFifo_3_29;
  wire       [5:0]    _zz_when_ArraySlice_l165_96;
  wire       [5:0]    _zz_when_ArraySlice_l165_96_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_96_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_96;
  wire       [6:0]    _zz_when_ArraySlice_l166_96_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_96_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_96_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_96_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_96_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_96;
  wire       [6:0]    _zz_when_ArraySlice_l113_96;
  wire       [6:0]    _zz_when_ArraySlice_l113_96_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_96_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_96_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_96_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_96;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_96_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_96_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_96_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_96;
  wire       [6:0]    _zz_when_ArraySlice_l118_96_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_96_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_96_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_96_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_96_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_96_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_96_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_96_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_96_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_97;
  wire       [5:0]    _zz_when_ArraySlice_l165_97_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_97_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_97;
  wire       [5:0]    _zz_when_ArraySlice_l166_97_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_97_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_97_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_97_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_97;
  wire       [6:0]    _zz_when_ArraySlice_l113_97;
  wire       [6:0]    _zz_when_ArraySlice_l113_97_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_97_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_97_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_97_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_97;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_97_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_97_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_97_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_97;
  wire       [6:0]    _zz_when_ArraySlice_l118_97_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_97_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_97_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_97_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_97_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_97_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_97_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_97_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_97_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_97_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_98;
  wire       [5:0]    _zz_when_ArraySlice_l165_98_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_98_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_98;
  wire       [5:0]    _zz_when_ArraySlice_l166_98_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_98_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_98_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_98_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_98;
  wire       [6:0]    _zz_when_ArraySlice_l113_98;
  wire       [6:0]    _zz_when_ArraySlice_l113_98_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_98_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_98_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_98_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_98;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_98_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_98_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_98_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_98;
  wire       [6:0]    _zz_when_ArraySlice_l118_98_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_98_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_98_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_98_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_98_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_98_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_98_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_98_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_98_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_98_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_99;
  wire       [5:0]    _zz_when_ArraySlice_l165_99_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_99_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_99;
  wire       [5:0]    _zz_when_ArraySlice_l166_99_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_99_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_99_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_99_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_99;
  wire       [6:0]    _zz_when_ArraySlice_l113_99;
  wire       [6:0]    _zz_when_ArraySlice_l113_99_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_99_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_99_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_99_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_99;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_99_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_99_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_99_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_99;
  wire       [6:0]    _zz_when_ArraySlice_l118_99_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_99_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_99_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_99_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_99_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_99_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_99_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_99_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_99_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_99_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_100;
  wire       [5:0]    _zz_when_ArraySlice_l165_100_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_100;
  wire       [5:0]    _zz_when_ArraySlice_l166_100_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_100_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_100_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_100;
  wire       [6:0]    _zz_when_ArraySlice_l113_100;
  wire       [6:0]    _zz_when_ArraySlice_l113_100_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_100_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_100_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_100_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_100;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_100_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_100_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_100_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_100;
  wire       [6:0]    _zz_when_ArraySlice_l118_100_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_100_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_100_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_100_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_100_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_100_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_100_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_100_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_100_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_101;
  wire       [5:0]    _zz_when_ArraySlice_l165_101_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_101;
  wire       [4:0]    _zz_when_ArraySlice_l166_101_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_101_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_101_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_101_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_101;
  wire       [6:0]    _zz_when_ArraySlice_l113_101;
  wire       [6:0]    _zz_when_ArraySlice_l113_101_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_101_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_101_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_101_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_101;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_101_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_101_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_101_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_101;
  wire       [6:0]    _zz_when_ArraySlice_l118_101_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_101_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_101_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_101_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_101_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_101_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_101_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_101_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_101_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_102;
  wire       [5:0]    _zz_when_ArraySlice_l165_102_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_102;
  wire       [4:0]    _zz_when_ArraySlice_l166_102_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_102_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_102_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_102_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_102;
  wire       [6:0]    _zz_when_ArraySlice_l113_102;
  wire       [6:0]    _zz_when_ArraySlice_l113_102_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_102_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_102_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_102_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_102;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_102_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_102_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_102_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_102;
  wire       [6:0]    _zz_when_ArraySlice_l118_102_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_102_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_102_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_102_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_102_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_102_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_102_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_102_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_102_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_103;
  wire       [5:0]    _zz_when_ArraySlice_l165_103_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_103;
  wire       [3:0]    _zz_when_ArraySlice_l166_103_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_103_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_103_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_103_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_103;
  wire       [6:0]    _zz_when_ArraySlice_l113_103;
  wire       [6:0]    _zz_when_ArraySlice_l113_103_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_103_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_103_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_103_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_103;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_103_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_103_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_103_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_103;
  wire       [6:0]    _zz_when_ArraySlice_l118_103_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_103_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_103_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_103_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_103_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_103_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_103_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_103_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_103_8;
  wire                _zz_when_ArraySlice_l444_3_1;
  wire                _zz_when_ArraySlice_l444_3_2;
  wire                _zz_when_ArraySlice_l444_3_3;
  wire                _zz_when_ArraySlice_l444_3_4;
  wire                _zz_when_ArraySlice_l444_3_5;
  wire                _zz_when_ArraySlice_l444_3_6;
  wire       [5:0]    _zz_selectReadFifo_3_30;
  wire       [0:0]    _zz_selectReadFifo_3_31;
  wire       [12:0]   _zz_when_ArraySlice_l448_3_1;
  wire       [12:0]   _zz_when_ArraySlice_l448_3_2;
  wire       [12:0]   _zz_when_ArraySlice_l448_3_3;
  wire       [0:0]    _zz_when_ArraySlice_l448_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l434_3;
  wire       [5:0]    _zz_when_ArraySlice_l434_3_1;
  wire       [4:0]    _zz_when_ArraySlice_l434_3_2;
  wire       [12:0]   _zz_when_ArraySlice_l455_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l455_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l455_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l455_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l455_3_5;
  wire       [5:0]    _zz_when_ArraySlice_l373_4;
  wire       [5:0]    _zz_when_ArraySlice_l373_4_1;
  reg        [6:0]    _zz_when_ArraySlice_l374_4;
  wire       [5:0]    _zz_when_ArraySlice_l374_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l374_4_2;
  wire       [5:0]    _zz__zz_outputStreamArrayData_4_valid;
  reg                 _zz_outputStreamArrayData_4_valid_2;
  reg        [31:0]   _zz_outputStreamArrayData_4_payload;
  wire       [6:0]    _zz_when_ArraySlice_l380_4_1;
  wire       [0:0]    _zz_when_ArraySlice_l380_4_2;
  reg        [6:0]    _zz_when_ArraySlice_l380_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l380_4_4;
  wire       [5:0]    _zz_when_ArraySlice_l380_4_5;
  wire       [12:0]   _zz_when_ArraySlice_l381_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l381_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l381_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l381_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l381_4_5;
  wire       [5:0]    _zz_selectReadFifo_4;
  wire       [5:0]    _zz_selectReadFifo_4_1;
  wire       [5:0]    _zz_selectReadFifo_4_2;
  wire       [0:0]    _zz_selectReadFifo_4_3;
  wire       [5:0]    _zz_selectReadFifo_4_4;
  wire       [0:0]    _zz_selectReadFifo_4_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_4;
  wire       [12:0]   _zz_when_ArraySlice_l384_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l384_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l384_4_3;
  reg        [6:0]    _zz_when_ArraySlice_l389_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l389_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l389_4_3;
  wire       [6:0]    _zz_when_ArraySlice_l389_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l389_4_5;
  wire       [12:0]   _zz_when_ArraySlice_l390_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l390_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l390_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l390_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l390_4_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_12;
  wire       [6:0]    _zz_when_ArraySlice_l95_12;
  wire       [6:0]    _zz_when_ArraySlice_l95_12_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_12_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_12_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_12_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_4_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_4_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_12;
  wire       [6:0]    _zz_when_ArraySlice_l99_12_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l392_4_3;
  wire       [6:0]    _zz_when_ArraySlice_l392_4_4;
  wire       [5:0]    _zz_selectReadFifo_4_6;
  wire       [5:0]    _zz_selectReadFifo_4_7;
  wire       [5:0]    _zz_selectReadFifo_4_8;
  wire       [0:0]    _zz_selectReadFifo_4_9;
  wire       [5:0]    _zz_selectReadFifo_4_10;
  wire       [5:0]    _zz_selectReadFifo_4_11;
  wire       [5:0]    _zz_selectReadFifo_4_12;
  wire       [0:0]    _zz_selectReadFifo_4_13;
  wire       [5:0]    _zz_when_ArraySlice_l165_104;
  wire       [5:0]    _zz_when_ArraySlice_l165_104_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_104_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_104;
  wire       [6:0]    _zz_when_ArraySlice_l166_104_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_104_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_104_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_104_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_104_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_104;
  wire       [6:0]    _zz_when_ArraySlice_l113_104;
  wire       [6:0]    _zz_when_ArraySlice_l113_104_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_104_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_104_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_104_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_104;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_104_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_104_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_104_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_104;
  wire       [6:0]    _zz_when_ArraySlice_l118_104_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_104_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_104_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_104_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_104_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_104_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_104_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_104_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_104_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_105;
  wire       [5:0]    _zz_when_ArraySlice_l165_105_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_105_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_105;
  wire       [5:0]    _zz_when_ArraySlice_l166_105_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_105_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_105_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_105_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_105;
  wire       [6:0]    _zz_when_ArraySlice_l113_105;
  wire       [6:0]    _zz_when_ArraySlice_l113_105_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_105_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_105_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_105_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_105;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_105_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_105_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_105_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_105;
  wire       [6:0]    _zz_when_ArraySlice_l118_105_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_105_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_105_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_105_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_105_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_105_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_105_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_105_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_105_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_105_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_106;
  wire       [5:0]    _zz_when_ArraySlice_l165_106_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_106_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_106;
  wire       [5:0]    _zz_when_ArraySlice_l166_106_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_106_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_106_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_106_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_106;
  wire       [6:0]    _zz_when_ArraySlice_l113_106;
  wire       [6:0]    _zz_when_ArraySlice_l113_106_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_106_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_106_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_106_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_106;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_106_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_106_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_106_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_106;
  wire       [6:0]    _zz_when_ArraySlice_l118_106_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_106_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_106_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_106_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_106_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_106_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_106_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_106_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_106_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_106_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_107;
  wire       [5:0]    _zz_when_ArraySlice_l165_107_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_107_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_107;
  wire       [5:0]    _zz_when_ArraySlice_l166_107_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_107_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_107_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_107_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_107;
  wire       [6:0]    _zz_when_ArraySlice_l113_107;
  wire       [6:0]    _zz_when_ArraySlice_l113_107_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_107_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_107_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_107_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_107;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_107_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_107_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_107_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_107;
  wire       [6:0]    _zz_when_ArraySlice_l118_107_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_107_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_107_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_107_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_107_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_107_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_107_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_107_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_107_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_107_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_108;
  wire       [5:0]    _zz_when_ArraySlice_l165_108_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_108;
  wire       [5:0]    _zz_when_ArraySlice_l166_108_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_108_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_108_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_108;
  wire       [6:0]    _zz_when_ArraySlice_l113_108;
  wire       [6:0]    _zz_when_ArraySlice_l113_108_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_108_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_108_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_108_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_108;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_108_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_108_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_108_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_108;
  wire       [6:0]    _zz_when_ArraySlice_l118_108_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_108_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_108_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_108_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_108_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_108_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_108_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_108_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_108_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_109;
  wire       [5:0]    _zz_when_ArraySlice_l165_109_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_109;
  wire       [4:0]    _zz_when_ArraySlice_l166_109_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_109_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_109_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_109_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_109;
  wire       [6:0]    _zz_when_ArraySlice_l113_109;
  wire       [6:0]    _zz_when_ArraySlice_l113_109_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_109_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_109_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_109_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_109;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_109_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_109_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_109_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_109;
  wire       [6:0]    _zz_when_ArraySlice_l118_109_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_109_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_109_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_109_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_109_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_109_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_109_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_109_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_109_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_110;
  wire       [5:0]    _zz_when_ArraySlice_l165_110_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_110;
  wire       [4:0]    _zz_when_ArraySlice_l166_110_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_110_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_110_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_110_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_110;
  wire       [6:0]    _zz_when_ArraySlice_l113_110;
  wire       [6:0]    _zz_when_ArraySlice_l113_110_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_110_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_110_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_110_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_110;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_110_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_110_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_110_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_110;
  wire       [6:0]    _zz_when_ArraySlice_l118_110_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_110_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_110_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_110_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_110_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_110_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_110_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_110_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_110_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_111;
  wire       [5:0]    _zz_when_ArraySlice_l165_111_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_111;
  wire       [3:0]    _zz_when_ArraySlice_l166_111_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_111_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_111_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_111_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_111;
  wire       [6:0]    _zz_when_ArraySlice_l113_111;
  wire       [6:0]    _zz_when_ArraySlice_l113_111_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_111_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_111_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_111_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_111;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_111_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_111_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_111_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_111;
  wire       [6:0]    _zz_when_ArraySlice_l118_111_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_111_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_111_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_111_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_111_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_111_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_111_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_111_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_111_8;
  wire                _zz_when_ArraySlice_l398_4_1;
  wire                _zz_when_ArraySlice_l398_4_2;
  wire                _zz_when_ArraySlice_l398_4_3;
  wire                _zz_when_ArraySlice_l398_4_4;
  wire                _zz_when_ArraySlice_l398_4_5;
  wire                _zz_when_ArraySlice_l398_4_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l401_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l401_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l401_4_4;
  wire       [5:0]    _zz_when_ArraySlice_l401_4_5;
  wire       [0:0]    _zz_when_ArraySlice_l401_4_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_4_7;
  wire       [5:0]    _zz_selectReadFifo_4_14;
  wire       [0:0]    _zz_selectReadFifo_4_15;
  wire       [12:0]   _zz_when_ArraySlice_l405_4;
  wire       [12:0]   _zz_when_ArraySlice_l405_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l405_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l405_4_3;
  reg        [6:0]    _zz_when_ArraySlice_l409_4;
  wire       [5:0]    _zz_when_ArraySlice_l409_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l409_4_2;
  wire       [12:0]   _zz_when_ArraySlice_l410_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l410_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l410_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l410_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l410_4_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_13;
  wire       [6:0]    _zz_when_ArraySlice_l95_13;
  wire       [6:0]    _zz_when_ArraySlice_l95_13_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_13_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_13_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_13_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_4_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_4_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_13;
  wire       [6:0]    _zz_when_ArraySlice_l99_13_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l412_4_3;
  wire       [6:0]    _zz_when_ArraySlice_l412_4_4;
  wire       [5:0]    _zz_selectReadFifo_4_16;
  wire       [5:0]    _zz_selectReadFifo_4_17;
  wire       [5:0]    _zz_selectReadFifo_4_18;
  wire       [0:0]    _zz_selectReadFifo_4_19;
  wire       [5:0]    _zz_selectReadFifo_4_20;
  wire       [5:0]    _zz_selectReadFifo_4_21;
  wire       [5:0]    _zz_selectReadFifo_4_22;
  wire       [0:0]    _zz_selectReadFifo_4_23;
  wire       [5:0]    _zz_when_ArraySlice_l165_112;
  wire       [5:0]    _zz_when_ArraySlice_l165_112_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_112_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_112;
  wire       [6:0]    _zz_when_ArraySlice_l166_112_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_112_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_112_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_112_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_112_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_112;
  wire       [6:0]    _zz_when_ArraySlice_l113_112;
  wire       [6:0]    _zz_when_ArraySlice_l113_112_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_112_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_112_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_112_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_112;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_112_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_112_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_112_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_112;
  wire       [6:0]    _zz_when_ArraySlice_l118_112_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_112_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_112_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_112_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_112_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_112_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_112_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_112_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_112_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_113;
  wire       [5:0]    _zz_when_ArraySlice_l165_113_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_113_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_113;
  wire       [5:0]    _zz_when_ArraySlice_l166_113_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_113_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_113_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_113_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_113;
  wire       [6:0]    _zz_when_ArraySlice_l113_113;
  wire       [6:0]    _zz_when_ArraySlice_l113_113_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_113_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_113_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_113_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_113;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_113_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_113_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_113_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_113;
  wire       [6:0]    _zz_when_ArraySlice_l118_113_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_113_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_113_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_113_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_113_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_113_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_113_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_113_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_113_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_113_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_114;
  wire       [5:0]    _zz_when_ArraySlice_l165_114_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_114_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_114;
  wire       [5:0]    _zz_when_ArraySlice_l166_114_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_114_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_114_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_114_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_114;
  wire       [6:0]    _zz_when_ArraySlice_l113_114;
  wire       [6:0]    _zz_when_ArraySlice_l113_114_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_114_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_114_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_114_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_114;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_114_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_114_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_114_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_114;
  wire       [6:0]    _zz_when_ArraySlice_l118_114_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_114_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_114_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_114_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_114_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_114_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_114_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_114_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_114_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_114_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_115;
  wire       [5:0]    _zz_when_ArraySlice_l165_115_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_115_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_115;
  wire       [5:0]    _zz_when_ArraySlice_l166_115_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_115_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_115_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_115_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_115;
  wire       [6:0]    _zz_when_ArraySlice_l113_115;
  wire       [6:0]    _zz_when_ArraySlice_l113_115_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_115_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_115_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_115_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_115;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_115_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_115_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_115_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_115;
  wire       [6:0]    _zz_when_ArraySlice_l118_115_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_115_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_115_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_115_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_115_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_115_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_115_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_115_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_115_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_115_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_116;
  wire       [5:0]    _zz_when_ArraySlice_l165_116_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_116;
  wire       [5:0]    _zz_when_ArraySlice_l166_116_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_116_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_116_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_116;
  wire       [6:0]    _zz_when_ArraySlice_l113_116;
  wire       [6:0]    _zz_when_ArraySlice_l113_116_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_116_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_116_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_116_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_116;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_116_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_116_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_116_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_116;
  wire       [6:0]    _zz_when_ArraySlice_l118_116_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_116_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_116_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_116_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_116_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_116_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_116_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_116_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_116_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_117;
  wire       [5:0]    _zz_when_ArraySlice_l165_117_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_117;
  wire       [4:0]    _zz_when_ArraySlice_l166_117_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_117_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_117_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_117_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_117;
  wire       [6:0]    _zz_when_ArraySlice_l113_117;
  wire       [6:0]    _zz_when_ArraySlice_l113_117_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_117_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_117_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_117_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_117;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_117_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_117_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_117_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_117;
  wire       [6:0]    _zz_when_ArraySlice_l118_117_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_117_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_117_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_117_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_117_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_117_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_117_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_117_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_117_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_118;
  wire       [5:0]    _zz_when_ArraySlice_l165_118_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_118;
  wire       [4:0]    _zz_when_ArraySlice_l166_118_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_118_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_118_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_118_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_118;
  wire       [6:0]    _zz_when_ArraySlice_l113_118;
  wire       [6:0]    _zz_when_ArraySlice_l113_118_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_118_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_118_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_118_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_118;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_118_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_118_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_118_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_118;
  wire       [6:0]    _zz_when_ArraySlice_l118_118_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_118_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_118_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_118_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_118_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_118_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_118_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_118_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_118_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_119;
  wire       [5:0]    _zz_when_ArraySlice_l165_119_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_119;
  wire       [3:0]    _zz_when_ArraySlice_l166_119_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_119_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_119_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_119_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_119;
  wire       [6:0]    _zz_when_ArraySlice_l113_119;
  wire       [6:0]    _zz_when_ArraySlice_l113_119_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_119_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_119_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_119_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_119;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_119_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_119_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_119_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_119;
  wire       [6:0]    _zz_when_ArraySlice_l118_119_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_119_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_119_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_119_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_119_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_119_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_119_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_119_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_119_8;
  wire                _zz_when_ArraySlice_l418_4_1;
  wire                _zz_when_ArraySlice_l418_4_2;
  wire                _zz_when_ArraySlice_l418_4_3;
  wire                _zz_when_ArraySlice_l418_4_4;
  wire                _zz_when_ArraySlice_l418_4_5;
  wire                _zz_when_ArraySlice_l418_4_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l421_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l421_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l421_4_4;
  wire       [5:0]    _zz_when_ArraySlice_l421_4_5;
  wire       [0:0]    _zz_when_ArraySlice_l421_4_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_4_7;
  wire       [5:0]    _zz_selectReadFifo_4_24;
  wire       [0:0]    _zz_selectReadFifo_4_25;
  wire       [12:0]   _zz_when_ArraySlice_l425_4;
  wire       [12:0]   _zz_when_ArraySlice_l425_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l425_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l425_4_3;
  wire       [12:0]   _zz_when_ArraySlice_l436_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l436_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l436_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l436_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l436_4_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_14;
  wire       [6:0]    _zz_when_ArraySlice_l95_14;
  wire       [6:0]    _zz_when_ArraySlice_l95_14_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_14_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_14_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_14_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_4_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_4_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_14;
  wire       [6:0]    _zz_when_ArraySlice_l99_14_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l437_4_3;
  wire       [6:0]    _zz_when_ArraySlice_l437_4_4;
  wire       [5:0]    _zz_selectReadFifo_4_26;
  wire       [5:0]    _zz_selectReadFifo_4_27;
  wire       [5:0]    _zz_selectReadFifo_4_28;
  wire       [0:0]    _zz_selectReadFifo_4_29;
  wire       [5:0]    _zz_when_ArraySlice_l165_120;
  wire       [5:0]    _zz_when_ArraySlice_l165_120_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_120_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_120;
  wire       [6:0]    _zz_when_ArraySlice_l166_120_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_120_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_120_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_120_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_120_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_120;
  wire       [6:0]    _zz_when_ArraySlice_l113_120;
  wire       [6:0]    _zz_when_ArraySlice_l113_120_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_120_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_120_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_120_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_120;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_120_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_120_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_120_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_120;
  wire       [6:0]    _zz_when_ArraySlice_l118_120_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_120_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_120_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_120_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_120_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_120_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_120_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_120_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_120_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_121;
  wire       [5:0]    _zz_when_ArraySlice_l165_121_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_121_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_121;
  wire       [5:0]    _zz_when_ArraySlice_l166_121_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_121_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_121_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_121_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_121;
  wire       [6:0]    _zz_when_ArraySlice_l113_121;
  wire       [6:0]    _zz_when_ArraySlice_l113_121_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_121_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_121_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_121_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_121;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_121_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_121_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_121_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_121;
  wire       [6:0]    _zz_when_ArraySlice_l118_121_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_121_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_121_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_121_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_121_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_121_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_121_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_121_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_121_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_121_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_122;
  wire       [5:0]    _zz_when_ArraySlice_l165_122_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_122_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_122;
  wire       [5:0]    _zz_when_ArraySlice_l166_122_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_122_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_122_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_122_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_122;
  wire       [6:0]    _zz_when_ArraySlice_l113_122;
  wire       [6:0]    _zz_when_ArraySlice_l113_122_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_122_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_122_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_122_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_122;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_122_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_122_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_122_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_122;
  wire       [6:0]    _zz_when_ArraySlice_l118_122_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_122_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_122_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_122_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_122_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_122_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_122_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_122_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_122_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_122_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_123;
  wire       [5:0]    _zz_when_ArraySlice_l165_123_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_123_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_123;
  wire       [5:0]    _zz_when_ArraySlice_l166_123_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_123_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_123_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_123_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_123;
  wire       [6:0]    _zz_when_ArraySlice_l113_123;
  wire       [6:0]    _zz_when_ArraySlice_l113_123_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_123_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_123_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_123_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_123;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_123_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_123_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_123_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_123;
  wire       [6:0]    _zz_when_ArraySlice_l118_123_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_123_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_123_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_123_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_123_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_123_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_123_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_123_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_123_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_123_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_124;
  wire       [5:0]    _zz_when_ArraySlice_l165_124_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_124;
  wire       [5:0]    _zz_when_ArraySlice_l166_124_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_124_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_124_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_124;
  wire       [6:0]    _zz_when_ArraySlice_l113_124;
  wire       [6:0]    _zz_when_ArraySlice_l113_124_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_124_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_124_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_124_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_124;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_124_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_124_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_124_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_124;
  wire       [6:0]    _zz_when_ArraySlice_l118_124_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_124_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_124_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_124_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_124_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_124_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_124_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_124_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_124_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_125;
  wire       [5:0]    _zz_when_ArraySlice_l165_125_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_125;
  wire       [4:0]    _zz_when_ArraySlice_l166_125_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_125_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_125_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_125_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_125;
  wire       [6:0]    _zz_when_ArraySlice_l113_125;
  wire       [6:0]    _zz_when_ArraySlice_l113_125_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_125_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_125_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_125_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_125;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_125_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_125_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_125_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_125;
  wire       [6:0]    _zz_when_ArraySlice_l118_125_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_125_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_125_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_125_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_125_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_125_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_125_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_125_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_125_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_126;
  wire       [5:0]    _zz_when_ArraySlice_l165_126_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_126;
  wire       [4:0]    _zz_when_ArraySlice_l166_126_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_126_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_126_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_126_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_126;
  wire       [6:0]    _zz_when_ArraySlice_l113_126;
  wire       [6:0]    _zz_when_ArraySlice_l113_126_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_126_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_126_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_126_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_126;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_126_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_126_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_126_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_126;
  wire       [6:0]    _zz_when_ArraySlice_l118_126_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_126_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_126_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_126_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_126_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_126_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_126_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_126_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_126_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_127;
  wire       [5:0]    _zz_when_ArraySlice_l165_127_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_127;
  wire       [3:0]    _zz_when_ArraySlice_l166_127_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_127_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_127_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_127_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_127;
  wire       [6:0]    _zz_when_ArraySlice_l113_127;
  wire       [6:0]    _zz_when_ArraySlice_l113_127_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_127_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_127_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_127_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_127;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_127_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_127_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_127_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_127;
  wire       [6:0]    _zz_when_ArraySlice_l118_127_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_127_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_127_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_127_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_127_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_127_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_127_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_127_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_127_8;
  wire                _zz_when_ArraySlice_l444_4_1;
  wire                _zz_when_ArraySlice_l444_4_2;
  wire                _zz_when_ArraySlice_l444_4_3;
  wire                _zz_when_ArraySlice_l444_4_4;
  wire                _zz_when_ArraySlice_l444_4_5;
  wire                _zz_when_ArraySlice_l444_4_6;
  wire       [5:0]    _zz_selectReadFifo_4_30;
  wire       [0:0]    _zz_selectReadFifo_4_31;
  wire       [12:0]   _zz_when_ArraySlice_l448_4;
  wire       [12:0]   _zz_when_ArraySlice_l448_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l448_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l448_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l434_4;
  wire       [5:0]    _zz_when_ArraySlice_l434_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l455_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l455_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l455_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l455_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l455_4_5;
  wire       [5:0]    _zz_when_ArraySlice_l373_5;
  wire       [5:0]    _zz_when_ArraySlice_l373_5_1;
  reg        [6:0]    _zz_when_ArraySlice_l374_5;
  wire       [5:0]    _zz_when_ArraySlice_l374_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l374_5_2;
  wire       [5:0]    _zz__zz_outputStreamArrayData_5_valid;
  reg                 _zz_outputStreamArrayData_5_valid_2;
  reg        [31:0]   _zz_outputStreamArrayData_5_payload;
  wire       [6:0]    _zz_when_ArraySlice_l380_5_1;
  wire       [0:0]    _zz_when_ArraySlice_l380_5_2;
  reg        [6:0]    _zz_when_ArraySlice_l380_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l380_5_4;
  wire       [5:0]    _zz_when_ArraySlice_l380_5_5;
  wire       [12:0]   _zz_when_ArraySlice_l381_5;
  wire       [5:0]    _zz_when_ArraySlice_l381_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l381_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l381_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l381_5_4;
  wire       [5:0]    _zz_selectReadFifo_5;
  wire       [5:0]    _zz_selectReadFifo_5_1;
  wire       [5:0]    _zz_selectReadFifo_5_2;
  wire       [0:0]    _zz_selectReadFifo_5_3;
  wire       [5:0]    _zz_selectReadFifo_5_4;
  wire       [0:0]    _zz_selectReadFifo_5_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l384_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l384_5_3;
  reg        [6:0]    _zz_when_ArraySlice_l389_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l389_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l389_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l389_5_4;
  wire       [0:0]    _zz_when_ArraySlice_l389_5_5;
  wire       [12:0]   _zz_when_ArraySlice_l390_5;
  wire       [5:0]    _zz_when_ArraySlice_l390_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l390_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l390_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l390_5_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_15;
  wire       [6:0]    _zz_when_ArraySlice_l95_15;
  wire       [6:0]    _zz_when_ArraySlice_l95_15_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_15_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_15_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_15_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_5_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_5_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_15;
  wire       [6:0]    _zz_when_ArraySlice_l99_15_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l392_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l392_5_4;
  wire       [5:0]    _zz_selectReadFifo_5_6;
  wire       [5:0]    _zz_selectReadFifo_5_7;
  wire       [5:0]    _zz_selectReadFifo_5_8;
  wire       [0:0]    _zz_selectReadFifo_5_9;
  wire       [5:0]    _zz_selectReadFifo_5_10;
  wire       [5:0]    _zz_selectReadFifo_5_11;
  wire       [5:0]    _zz_selectReadFifo_5_12;
  wire       [0:0]    _zz_selectReadFifo_5_13;
  wire       [5:0]    _zz_when_ArraySlice_l165_128;
  wire       [5:0]    _zz_when_ArraySlice_l165_128_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_128_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_128;
  wire       [6:0]    _zz_when_ArraySlice_l166_128_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_128_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_128_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_128_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_128_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_128;
  wire       [6:0]    _zz_when_ArraySlice_l113_128;
  wire       [6:0]    _zz_when_ArraySlice_l113_128_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_128_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_128_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_128_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_128;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_128_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_128_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_128_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_128;
  wire       [6:0]    _zz_when_ArraySlice_l118_128_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_128_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_128_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_128_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_128_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_128_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_128_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_128_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_128_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_129;
  wire       [5:0]    _zz_when_ArraySlice_l165_129_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_129_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_129;
  wire       [5:0]    _zz_when_ArraySlice_l166_129_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_129_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_129_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_129_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_129;
  wire       [6:0]    _zz_when_ArraySlice_l113_129;
  wire       [6:0]    _zz_when_ArraySlice_l113_129_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_129_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_129_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_129_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_129;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_129_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_129_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_129_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_129;
  wire       [6:0]    _zz_when_ArraySlice_l118_129_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_129_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_129_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_129_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_129_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_129_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_129_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_129_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_129_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_129_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_130;
  wire       [5:0]    _zz_when_ArraySlice_l165_130_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_130_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_130;
  wire       [5:0]    _zz_when_ArraySlice_l166_130_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_130_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_130_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_130_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_130;
  wire       [6:0]    _zz_when_ArraySlice_l113_130;
  wire       [6:0]    _zz_when_ArraySlice_l113_130_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_130_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_130_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_130_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_130;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_130_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_130_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_130_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_130;
  wire       [6:0]    _zz_when_ArraySlice_l118_130_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_130_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_130_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_130_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_130_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_130_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_130_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_130_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_130_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_130_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_131;
  wire       [5:0]    _zz_when_ArraySlice_l165_131_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_131_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_131;
  wire       [5:0]    _zz_when_ArraySlice_l166_131_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_131_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_131_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_131_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_131;
  wire       [6:0]    _zz_when_ArraySlice_l113_131;
  wire       [6:0]    _zz_when_ArraySlice_l113_131_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_131_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_131_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_131_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_131;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_131_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_131_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_131_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_131;
  wire       [6:0]    _zz_when_ArraySlice_l118_131_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_131_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_131_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_131_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_131_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_131_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_131_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_131_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_131_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_131_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_132;
  wire       [5:0]    _zz_when_ArraySlice_l165_132_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_132;
  wire       [5:0]    _zz_when_ArraySlice_l166_132_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_132_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_132_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_132;
  wire       [6:0]    _zz_when_ArraySlice_l113_132;
  wire       [6:0]    _zz_when_ArraySlice_l113_132_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_132_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_132_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_132_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_132;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_132_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_132_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_132_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_132;
  wire       [6:0]    _zz_when_ArraySlice_l118_132_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_132_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_132_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_132_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_132_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_132_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_132_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_132_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_132_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_133;
  wire       [5:0]    _zz_when_ArraySlice_l165_133_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_133;
  wire       [4:0]    _zz_when_ArraySlice_l166_133_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_133_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_133_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_133_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_133;
  wire       [6:0]    _zz_when_ArraySlice_l113_133;
  wire       [6:0]    _zz_when_ArraySlice_l113_133_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_133_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_133_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_133_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_133;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_133_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_133_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_133_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_133;
  wire       [6:0]    _zz_when_ArraySlice_l118_133_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_133_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_133_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_133_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_133_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_133_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_133_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_133_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_133_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_134;
  wire       [5:0]    _zz_when_ArraySlice_l165_134_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_134;
  wire       [4:0]    _zz_when_ArraySlice_l166_134_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_134_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_134_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_134_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_134;
  wire       [6:0]    _zz_when_ArraySlice_l113_134;
  wire       [6:0]    _zz_when_ArraySlice_l113_134_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_134_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_134_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_134_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_134;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_134_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_134_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_134_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_134;
  wire       [6:0]    _zz_when_ArraySlice_l118_134_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_134_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_134_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_134_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_134_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_134_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_134_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_134_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_134_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_135;
  wire       [5:0]    _zz_when_ArraySlice_l165_135_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_135;
  wire       [3:0]    _zz_when_ArraySlice_l166_135_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_135_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_135_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_135_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_135;
  wire       [6:0]    _zz_when_ArraySlice_l113_135;
  wire       [6:0]    _zz_when_ArraySlice_l113_135_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_135_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_135_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_135_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_135;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_135_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_135_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_135_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_135;
  wire       [6:0]    _zz_when_ArraySlice_l118_135_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_135_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_135_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_135_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_135_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_135_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_135_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_135_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_135_8;
  wire                _zz_when_ArraySlice_l398_5_1;
  wire                _zz_when_ArraySlice_l398_5_2;
  wire                _zz_when_ArraySlice_l398_5_3;
  wire                _zz_when_ArraySlice_l398_5_4;
  wire                _zz_when_ArraySlice_l398_5_5;
  wire                _zz_when_ArraySlice_l398_5_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l401_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l401_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l401_5_4;
  wire       [5:0]    _zz_when_ArraySlice_l401_5_5;
  wire       [0:0]    _zz_when_ArraySlice_l401_5_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_5_7;
  wire       [5:0]    _zz_selectReadFifo_5_14;
  wire       [0:0]    _zz_selectReadFifo_5_15;
  wire       [12:0]   _zz_when_ArraySlice_l405_5;
  wire       [12:0]   _zz_when_ArraySlice_l405_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l405_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l405_5_3;
  reg        [6:0]    _zz_when_ArraySlice_l409_5;
  wire       [5:0]    _zz_when_ArraySlice_l409_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l409_5_2;
  wire       [12:0]   _zz_when_ArraySlice_l410_5;
  wire       [5:0]    _zz_when_ArraySlice_l410_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l410_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l410_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l410_5_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_16;
  wire       [6:0]    _zz_when_ArraySlice_l95_16;
  wire       [6:0]    _zz_when_ArraySlice_l95_16_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_16_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_16_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_16_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_5_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_5_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_16;
  wire       [6:0]    _zz_when_ArraySlice_l99_16_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l412_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l412_5_4;
  wire       [5:0]    _zz_selectReadFifo_5_16;
  wire       [5:0]    _zz_selectReadFifo_5_17;
  wire       [5:0]    _zz_selectReadFifo_5_18;
  wire       [0:0]    _zz_selectReadFifo_5_19;
  wire       [5:0]    _zz_selectReadFifo_5_20;
  wire       [5:0]    _zz_selectReadFifo_5_21;
  wire       [5:0]    _zz_selectReadFifo_5_22;
  wire       [0:0]    _zz_selectReadFifo_5_23;
  wire       [5:0]    _zz_when_ArraySlice_l165_136;
  wire       [5:0]    _zz_when_ArraySlice_l165_136_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_136_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_136;
  wire       [6:0]    _zz_when_ArraySlice_l166_136_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_136_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_136_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_136_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_136_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_136;
  wire       [6:0]    _zz_when_ArraySlice_l113_136;
  wire       [6:0]    _zz_when_ArraySlice_l113_136_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_136_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_136_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_136_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_136;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_136_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_136_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_136_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_136;
  wire       [6:0]    _zz_when_ArraySlice_l118_136_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_136_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_136_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_136_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_136_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_136_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_136_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_136_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_136_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_137;
  wire       [5:0]    _zz_when_ArraySlice_l165_137_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_137_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_137;
  wire       [5:0]    _zz_when_ArraySlice_l166_137_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_137_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_137_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_137_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_137;
  wire       [6:0]    _zz_when_ArraySlice_l113_137;
  wire       [6:0]    _zz_when_ArraySlice_l113_137_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_137_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_137_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_137_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_137;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_137_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_137_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_137_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_137;
  wire       [6:0]    _zz_when_ArraySlice_l118_137_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_137_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_137_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_137_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_137_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_137_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_137_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_137_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_137_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_137_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_138;
  wire       [5:0]    _zz_when_ArraySlice_l165_138_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_138_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_138;
  wire       [5:0]    _zz_when_ArraySlice_l166_138_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_138_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_138_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_138_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_138;
  wire       [6:0]    _zz_when_ArraySlice_l113_138;
  wire       [6:0]    _zz_when_ArraySlice_l113_138_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_138_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_138_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_138_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_138;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_138_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_138_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_138_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_138;
  wire       [6:0]    _zz_when_ArraySlice_l118_138_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_138_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_138_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_138_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_138_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_138_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_138_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_138_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_138_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_138_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_139;
  wire       [5:0]    _zz_when_ArraySlice_l165_139_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_139_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_139;
  wire       [5:0]    _zz_when_ArraySlice_l166_139_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_139_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_139_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_139_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_139;
  wire       [6:0]    _zz_when_ArraySlice_l113_139;
  wire       [6:0]    _zz_when_ArraySlice_l113_139_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_139_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_139_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_139_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_139;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_139_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_139_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_139_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_139;
  wire       [6:0]    _zz_when_ArraySlice_l118_139_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_139_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_139_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_139_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_139_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_139_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_139_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_139_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_139_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_139_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_140;
  wire       [5:0]    _zz_when_ArraySlice_l165_140_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_140;
  wire       [5:0]    _zz_when_ArraySlice_l166_140_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_140_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_140_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_140;
  wire       [6:0]    _zz_when_ArraySlice_l113_140;
  wire       [6:0]    _zz_when_ArraySlice_l113_140_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_140_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_140_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_140_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_140;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_140_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_140_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_140_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_140;
  wire       [6:0]    _zz_when_ArraySlice_l118_140_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_140_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_140_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_140_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_140_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_140_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_140_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_140_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_140_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_141;
  wire       [5:0]    _zz_when_ArraySlice_l165_141_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_141;
  wire       [4:0]    _zz_when_ArraySlice_l166_141_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_141_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_141_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_141_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_141;
  wire       [6:0]    _zz_when_ArraySlice_l113_141;
  wire       [6:0]    _zz_when_ArraySlice_l113_141_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_141_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_141_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_141_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_141;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_141_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_141_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_141_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_141;
  wire       [6:0]    _zz_when_ArraySlice_l118_141_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_141_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_141_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_141_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_141_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_141_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_141_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_141_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_141_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_142;
  wire       [5:0]    _zz_when_ArraySlice_l165_142_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_142;
  wire       [4:0]    _zz_when_ArraySlice_l166_142_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_142_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_142_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_142_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_142;
  wire       [6:0]    _zz_when_ArraySlice_l113_142;
  wire       [6:0]    _zz_when_ArraySlice_l113_142_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_142_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_142_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_142_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_142;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_142_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_142_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_142_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_142;
  wire       [6:0]    _zz_when_ArraySlice_l118_142_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_142_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_142_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_142_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_142_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_142_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_142_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_142_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_142_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_143;
  wire       [5:0]    _zz_when_ArraySlice_l165_143_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_143;
  wire       [3:0]    _zz_when_ArraySlice_l166_143_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_143_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_143_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_143_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_143;
  wire       [6:0]    _zz_when_ArraySlice_l113_143;
  wire       [6:0]    _zz_when_ArraySlice_l113_143_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_143_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_143_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_143_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_143;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_143_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_143_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_143_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_143;
  wire       [6:0]    _zz_when_ArraySlice_l118_143_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_143_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_143_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_143_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_143_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_143_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_143_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_143_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_143_8;
  wire                _zz_when_ArraySlice_l418_5_1;
  wire                _zz_when_ArraySlice_l418_5_2;
  wire                _zz_when_ArraySlice_l418_5_3;
  wire                _zz_when_ArraySlice_l418_5_4;
  wire                _zz_when_ArraySlice_l418_5_5;
  wire                _zz_when_ArraySlice_l418_5_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l421_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l421_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l421_5_4;
  wire       [5:0]    _zz_when_ArraySlice_l421_5_5;
  wire       [0:0]    _zz_when_ArraySlice_l421_5_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_5_7;
  wire       [5:0]    _zz_selectReadFifo_5_24;
  wire       [0:0]    _zz_selectReadFifo_5_25;
  wire       [12:0]   _zz_when_ArraySlice_l425_5;
  wire       [12:0]   _zz_when_ArraySlice_l425_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l425_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l425_5_3;
  wire       [12:0]   _zz_when_ArraySlice_l436_5;
  wire       [5:0]    _zz_when_ArraySlice_l436_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l436_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l436_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l436_5_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_17;
  wire       [6:0]    _zz_when_ArraySlice_l95_17;
  wire       [6:0]    _zz_when_ArraySlice_l95_17_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_17_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_17_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_17_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_5_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_5_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_17;
  wire       [6:0]    _zz_when_ArraySlice_l99_17_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l437_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l437_5_4;
  wire       [5:0]    _zz_selectReadFifo_5_26;
  wire       [5:0]    _zz_selectReadFifo_5_27;
  wire       [5:0]    _zz_selectReadFifo_5_28;
  wire       [0:0]    _zz_selectReadFifo_5_29;
  wire       [5:0]    _zz_when_ArraySlice_l165_144;
  wire       [5:0]    _zz_when_ArraySlice_l165_144_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_144_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_144;
  wire       [6:0]    _zz_when_ArraySlice_l166_144_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_144_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_144_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_144_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_144_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_144;
  wire       [6:0]    _zz_when_ArraySlice_l113_144;
  wire       [6:0]    _zz_when_ArraySlice_l113_144_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_144_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_144_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_144_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_144;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_144_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_144_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_144_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_144;
  wire       [6:0]    _zz_when_ArraySlice_l118_144_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_144_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_144_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_144_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_144_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_144_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_144_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_144_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_144_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_145;
  wire       [5:0]    _zz_when_ArraySlice_l165_145_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_145_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_145;
  wire       [5:0]    _zz_when_ArraySlice_l166_145_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_145_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_145_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_145_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_145;
  wire       [6:0]    _zz_when_ArraySlice_l113_145;
  wire       [6:0]    _zz_when_ArraySlice_l113_145_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_145_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_145_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_145_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_145;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_145_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_145_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_145_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_145;
  wire       [6:0]    _zz_when_ArraySlice_l118_145_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_145_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_145_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_145_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_145_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_145_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_145_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_145_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_145_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_145_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_146;
  wire       [5:0]    _zz_when_ArraySlice_l165_146_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_146_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_146;
  wire       [5:0]    _zz_when_ArraySlice_l166_146_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_146_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_146_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_146_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_146;
  wire       [6:0]    _zz_when_ArraySlice_l113_146;
  wire       [6:0]    _zz_when_ArraySlice_l113_146_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_146_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_146_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_146_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_146;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_146_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_146_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_146_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_146;
  wire       [6:0]    _zz_when_ArraySlice_l118_146_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_146_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_146_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_146_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_146_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_146_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_146_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_146_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_146_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_146_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_147;
  wire       [5:0]    _zz_when_ArraySlice_l165_147_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_147_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_147;
  wire       [5:0]    _zz_when_ArraySlice_l166_147_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_147_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_147_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_147_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_147;
  wire       [6:0]    _zz_when_ArraySlice_l113_147;
  wire       [6:0]    _zz_when_ArraySlice_l113_147_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_147_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_147_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_147_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_147;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_147_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_147_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_147_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_147;
  wire       [6:0]    _zz_when_ArraySlice_l118_147_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_147_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_147_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_147_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_147_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_147_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_147_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_147_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_147_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_147_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_148;
  wire       [5:0]    _zz_when_ArraySlice_l165_148_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_148;
  wire       [5:0]    _zz_when_ArraySlice_l166_148_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_148_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_148_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_148;
  wire       [6:0]    _zz_when_ArraySlice_l113_148;
  wire       [6:0]    _zz_when_ArraySlice_l113_148_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_148_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_148_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_148_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_148;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_148_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_148_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_148_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_148;
  wire       [6:0]    _zz_when_ArraySlice_l118_148_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_148_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_148_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_148_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_148_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_148_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_148_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_148_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_148_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_149;
  wire       [5:0]    _zz_when_ArraySlice_l165_149_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_149;
  wire       [4:0]    _zz_when_ArraySlice_l166_149_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_149_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_149_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_149_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_149;
  wire       [6:0]    _zz_when_ArraySlice_l113_149;
  wire       [6:0]    _zz_when_ArraySlice_l113_149_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_149_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_149_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_149_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_149;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_149_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_149_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_149_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_149;
  wire       [6:0]    _zz_when_ArraySlice_l118_149_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_149_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_149_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_149_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_149_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_149_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_149_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_149_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_149_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_150;
  wire       [5:0]    _zz_when_ArraySlice_l165_150_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_150;
  wire       [4:0]    _zz_when_ArraySlice_l166_150_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_150_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_150_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_150_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_150;
  wire       [6:0]    _zz_when_ArraySlice_l113_150;
  wire       [6:0]    _zz_when_ArraySlice_l113_150_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_150_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_150_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_150_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_150;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_150_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_150_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_150_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_150;
  wire       [6:0]    _zz_when_ArraySlice_l118_150_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_150_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_150_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_150_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_150_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_150_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_150_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_150_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_150_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_151;
  wire       [5:0]    _zz_when_ArraySlice_l165_151_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_151;
  wire       [3:0]    _zz_when_ArraySlice_l166_151_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_151_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_151_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_151_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_151;
  wire       [6:0]    _zz_when_ArraySlice_l113_151;
  wire       [6:0]    _zz_when_ArraySlice_l113_151_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_151_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_151_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_151_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_151;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_151_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_151_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_151_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_151;
  wire       [6:0]    _zz_when_ArraySlice_l118_151_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_151_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_151_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_151_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_151_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_151_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_151_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_151_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_151_8;
  wire                _zz_when_ArraySlice_l444_5_1;
  wire                _zz_when_ArraySlice_l444_5_2;
  wire                _zz_when_ArraySlice_l444_5_3;
  wire                _zz_when_ArraySlice_l444_5_4;
  wire                _zz_when_ArraySlice_l444_5_5;
  wire                _zz_when_ArraySlice_l444_5_6;
  wire       [5:0]    _zz_selectReadFifo_5_30;
  wire       [0:0]    _zz_selectReadFifo_5_31;
  wire       [12:0]   _zz_when_ArraySlice_l448_5;
  wire       [12:0]   _zz_when_ArraySlice_l448_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l448_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l448_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l434_5;
  wire       [5:0]    _zz_when_ArraySlice_l434_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l455_5;
  wire       [5:0]    _zz_when_ArraySlice_l455_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l455_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l455_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l455_5_4;
  wire       [5:0]    _zz_when_ArraySlice_l373_6;
  wire       [5:0]    _zz_when_ArraySlice_l373_6_1;
  reg        [6:0]    _zz_when_ArraySlice_l374_6;
  wire       [5:0]    _zz_when_ArraySlice_l374_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l374_6_2;
  wire       [5:0]    _zz__zz_outputStreamArrayData_6_valid;
  reg                 _zz_outputStreamArrayData_6_valid_2;
  reg        [31:0]   _zz_outputStreamArrayData_6_payload;
  wire       [6:0]    _zz_when_ArraySlice_l380_6;
  wire       [0:0]    _zz_when_ArraySlice_l380_6_1;
  reg        [6:0]    _zz_when_ArraySlice_l380_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l380_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l380_6_4;
  wire       [12:0]   _zz_when_ArraySlice_l381_6;
  wire       [5:0]    _zz_when_ArraySlice_l381_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l381_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l381_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l381_6_4;
  wire       [5:0]    _zz_selectReadFifo_6;
  wire       [5:0]    _zz_selectReadFifo_6_1;
  wire       [5:0]    _zz_selectReadFifo_6_2;
  wire       [0:0]    _zz_selectReadFifo_6_3;
  wire       [5:0]    _zz_selectReadFifo_6_4;
  wire       [0:0]    _zz_selectReadFifo_6_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_6;
  wire       [12:0]   _zz_when_ArraySlice_l384_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l384_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l384_6_3;
  reg        [6:0]    _zz_when_ArraySlice_l389_6;
  wire       [5:0]    _zz_when_ArraySlice_l389_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l389_6_2;
  wire       [6:0]    _zz_when_ArraySlice_l389_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l389_6_4;
  wire       [12:0]   _zz_when_ArraySlice_l390_6;
  wire       [5:0]    _zz_when_ArraySlice_l390_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l390_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l390_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l390_6_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_18;
  wire       [6:0]    _zz_when_ArraySlice_l95_18;
  wire       [6:0]    _zz_when_ArraySlice_l95_18_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_18_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_18_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_18_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_6;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_6_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_6_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_18;
  wire       [6:0]    _zz_when_ArraySlice_l99_18_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l392_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l392_6_4;
  wire       [5:0]    _zz_selectReadFifo_6_6;
  wire       [5:0]    _zz_selectReadFifo_6_7;
  wire       [5:0]    _zz_selectReadFifo_6_8;
  wire       [0:0]    _zz_selectReadFifo_6_9;
  wire       [5:0]    _zz_selectReadFifo_6_10;
  wire       [5:0]    _zz_selectReadFifo_6_11;
  wire       [5:0]    _zz_selectReadFifo_6_12;
  wire       [0:0]    _zz_selectReadFifo_6_13;
  wire       [5:0]    _zz_when_ArraySlice_l165_152;
  wire       [5:0]    _zz_when_ArraySlice_l165_152_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_152_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_152;
  wire       [6:0]    _zz_when_ArraySlice_l166_152_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_152_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_152_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_152_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_152_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_152;
  wire       [6:0]    _zz_when_ArraySlice_l113_152;
  wire       [6:0]    _zz_when_ArraySlice_l113_152_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_152_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_152_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_152_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_152;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_152_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_152_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_152_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_152;
  wire       [6:0]    _zz_when_ArraySlice_l118_152_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_152_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_152_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_152_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_152_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_152_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_152_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_152_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_152_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_153;
  wire       [5:0]    _zz_when_ArraySlice_l165_153_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_153_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_153;
  wire       [5:0]    _zz_when_ArraySlice_l166_153_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_153_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_153_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_153_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_153;
  wire       [6:0]    _zz_when_ArraySlice_l113_153;
  wire       [6:0]    _zz_when_ArraySlice_l113_153_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_153_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_153_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_153_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_153;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_153_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_153_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_153_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_153;
  wire       [6:0]    _zz_when_ArraySlice_l118_153_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_153_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_153_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_153_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_153_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_153_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_153_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_153_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_153_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_153_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_154;
  wire       [5:0]    _zz_when_ArraySlice_l165_154_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_154_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_154;
  wire       [5:0]    _zz_when_ArraySlice_l166_154_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_154_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_154_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_154_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_154;
  wire       [6:0]    _zz_when_ArraySlice_l113_154;
  wire       [6:0]    _zz_when_ArraySlice_l113_154_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_154_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_154_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_154_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_154;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_154_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_154_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_154_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_154;
  wire       [6:0]    _zz_when_ArraySlice_l118_154_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_154_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_154_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_154_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_154_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_154_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_154_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_154_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_154_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_154_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_155;
  wire       [5:0]    _zz_when_ArraySlice_l165_155_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_155_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_155;
  wire       [5:0]    _zz_when_ArraySlice_l166_155_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_155_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_155_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_155_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_155;
  wire       [6:0]    _zz_when_ArraySlice_l113_155;
  wire       [6:0]    _zz_when_ArraySlice_l113_155_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_155_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_155_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_155_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_155;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_155_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_155_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_155_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_155;
  wire       [6:0]    _zz_when_ArraySlice_l118_155_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_155_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_155_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_155_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_155_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_155_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_155_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_155_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_155_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_155_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_156;
  wire       [5:0]    _zz_when_ArraySlice_l165_156_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_156;
  wire       [5:0]    _zz_when_ArraySlice_l166_156_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_156_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_156_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_156;
  wire       [6:0]    _zz_when_ArraySlice_l113_156;
  wire       [6:0]    _zz_when_ArraySlice_l113_156_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_156_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_156_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_156_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_156;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_156_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_156_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_156_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_156;
  wire       [6:0]    _zz_when_ArraySlice_l118_156_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_156_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_156_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_156_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_156_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_156_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_156_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_156_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_156_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_157;
  wire       [5:0]    _zz_when_ArraySlice_l165_157_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_157;
  wire       [4:0]    _zz_when_ArraySlice_l166_157_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_157_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_157_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_157_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_157;
  wire       [6:0]    _zz_when_ArraySlice_l113_157;
  wire       [6:0]    _zz_when_ArraySlice_l113_157_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_157_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_157_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_157_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_157;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_157_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_157_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_157_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_157;
  wire       [6:0]    _zz_when_ArraySlice_l118_157_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_157_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_157_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_157_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_157_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_157_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_157_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_157_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_157_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_158;
  wire       [5:0]    _zz_when_ArraySlice_l165_158_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_158;
  wire       [4:0]    _zz_when_ArraySlice_l166_158_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_158_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_158_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_158_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_158;
  wire       [6:0]    _zz_when_ArraySlice_l113_158;
  wire       [6:0]    _zz_when_ArraySlice_l113_158_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_158_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_158_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_158_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_158;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_158_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_158_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_158_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_158;
  wire       [6:0]    _zz_when_ArraySlice_l118_158_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_158_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_158_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_158_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_158_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_158_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_158_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_158_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_158_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_159;
  wire       [5:0]    _zz_when_ArraySlice_l165_159_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_159;
  wire       [3:0]    _zz_when_ArraySlice_l166_159_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_159_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_159_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_159_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_159;
  wire       [6:0]    _zz_when_ArraySlice_l113_159;
  wire       [6:0]    _zz_when_ArraySlice_l113_159_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_159_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_159_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_159_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_159;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_159_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_159_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_159_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_159;
  wire       [6:0]    _zz_when_ArraySlice_l118_159_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_159_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_159_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_159_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_159_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_159_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_159_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_159_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_159_8;
  wire                _zz_when_ArraySlice_l398_6_1;
  wire                _zz_when_ArraySlice_l398_6_2;
  wire                _zz_when_ArraySlice_l398_6_3;
  wire                _zz_when_ArraySlice_l398_6_4;
  wire                _zz_when_ArraySlice_l398_6_5;
  wire                _zz_when_ArraySlice_l398_6_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l401_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l401_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l401_6_4;
  wire       [5:0]    _zz_when_ArraySlice_l401_6_5;
  wire       [0:0]    _zz_when_ArraySlice_l401_6_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_6_7;
  wire       [5:0]    _zz_selectReadFifo_6_14;
  wire       [0:0]    _zz_selectReadFifo_6_15;
  wire       [12:0]   _zz_when_ArraySlice_l405_6;
  wire       [12:0]   _zz_when_ArraySlice_l405_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l405_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l405_6_3;
  reg        [6:0]    _zz_when_ArraySlice_l409_6;
  wire       [5:0]    _zz_when_ArraySlice_l409_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l409_6_2;
  wire       [12:0]   _zz_when_ArraySlice_l410_6;
  wire       [5:0]    _zz_when_ArraySlice_l410_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l410_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l410_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l410_6_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_19;
  wire       [6:0]    _zz_when_ArraySlice_l95_19;
  wire       [6:0]    _zz_when_ArraySlice_l95_19_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_19_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_19_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_19_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_6;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_6_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_6_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_19;
  wire       [6:0]    _zz_when_ArraySlice_l99_19_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l412_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l412_6_4;
  wire       [5:0]    _zz_selectReadFifo_6_16;
  wire       [5:0]    _zz_selectReadFifo_6_17;
  wire       [5:0]    _zz_selectReadFifo_6_18;
  wire       [0:0]    _zz_selectReadFifo_6_19;
  wire       [5:0]    _zz_selectReadFifo_6_20;
  wire       [5:0]    _zz_selectReadFifo_6_21;
  wire       [5:0]    _zz_selectReadFifo_6_22;
  wire       [0:0]    _zz_selectReadFifo_6_23;
  wire       [5:0]    _zz_when_ArraySlice_l165_160;
  wire       [5:0]    _zz_when_ArraySlice_l165_160_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_160_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_160;
  wire       [6:0]    _zz_when_ArraySlice_l166_160_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_160_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_160_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_160_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_160_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_160;
  wire       [6:0]    _zz_when_ArraySlice_l113_160;
  wire       [6:0]    _zz_when_ArraySlice_l113_160_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_160_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_160_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_160_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_160;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_160_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_160_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_160_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_160;
  wire       [6:0]    _zz_when_ArraySlice_l118_160_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_160_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_160_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_160_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_160_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_160_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_160_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_160_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_160_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_161;
  wire       [5:0]    _zz_when_ArraySlice_l165_161_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_161_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_161;
  wire       [5:0]    _zz_when_ArraySlice_l166_161_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_161_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_161_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_161_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_161;
  wire       [6:0]    _zz_when_ArraySlice_l113_161;
  wire       [6:0]    _zz_when_ArraySlice_l113_161_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_161_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_161_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_161_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_161;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_161_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_161_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_161_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_161;
  wire       [6:0]    _zz_when_ArraySlice_l118_161_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_161_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_161_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_161_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_161_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_161_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_161_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_161_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_161_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_161_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_162;
  wire       [5:0]    _zz_when_ArraySlice_l165_162_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_162_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_162;
  wire       [5:0]    _zz_when_ArraySlice_l166_162_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_162_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_162_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_162_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_162;
  wire       [6:0]    _zz_when_ArraySlice_l113_162;
  wire       [6:0]    _zz_when_ArraySlice_l113_162_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_162_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_162_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_162_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_162;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_162_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_162_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_162_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_162;
  wire       [6:0]    _zz_when_ArraySlice_l118_162_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_162_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_162_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_162_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_162_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_162_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_162_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_162_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_162_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_162_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_163;
  wire       [5:0]    _zz_when_ArraySlice_l165_163_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_163_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_163;
  wire       [5:0]    _zz_when_ArraySlice_l166_163_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_163_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_163_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_163_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_163;
  wire       [6:0]    _zz_when_ArraySlice_l113_163;
  wire       [6:0]    _zz_when_ArraySlice_l113_163_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_163_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_163_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_163_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_163;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_163_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_163_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_163_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_163;
  wire       [6:0]    _zz_when_ArraySlice_l118_163_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_163_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_163_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_163_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_163_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_163_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_163_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_163_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_163_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_163_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_164;
  wire       [5:0]    _zz_when_ArraySlice_l165_164_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_164;
  wire       [5:0]    _zz_when_ArraySlice_l166_164_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_164_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_164_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_164;
  wire       [6:0]    _zz_when_ArraySlice_l113_164;
  wire       [6:0]    _zz_when_ArraySlice_l113_164_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_164_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_164_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_164_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_164;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_164_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_164_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_164_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_164;
  wire       [6:0]    _zz_when_ArraySlice_l118_164_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_164_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_164_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_164_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_164_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_164_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_164_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_164_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_164_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_165;
  wire       [5:0]    _zz_when_ArraySlice_l165_165_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_165;
  wire       [4:0]    _zz_when_ArraySlice_l166_165_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_165_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_165_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_165_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_165;
  wire       [6:0]    _zz_when_ArraySlice_l113_165;
  wire       [6:0]    _zz_when_ArraySlice_l113_165_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_165_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_165_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_165_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_165;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_165_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_165_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_165_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_165;
  wire       [6:0]    _zz_when_ArraySlice_l118_165_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_165_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_165_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_165_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_165_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_165_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_165_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_165_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_165_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_166;
  wire       [5:0]    _zz_when_ArraySlice_l165_166_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_166;
  wire       [4:0]    _zz_when_ArraySlice_l166_166_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_166_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_166_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_166_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_166;
  wire       [6:0]    _zz_when_ArraySlice_l113_166;
  wire       [6:0]    _zz_when_ArraySlice_l113_166_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_166_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_166_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_166_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_166;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_166_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_166_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_166_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_166;
  wire       [6:0]    _zz_when_ArraySlice_l118_166_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_166_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_166_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_166_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_166_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_166_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_166_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_166_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_166_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_167;
  wire       [5:0]    _zz_when_ArraySlice_l165_167_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_167;
  wire       [3:0]    _zz_when_ArraySlice_l166_167_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_167_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_167_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_167_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_167;
  wire       [6:0]    _zz_when_ArraySlice_l113_167;
  wire       [6:0]    _zz_when_ArraySlice_l113_167_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_167_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_167_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_167_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_167;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_167_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_167_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_167_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_167;
  wire       [6:0]    _zz_when_ArraySlice_l118_167_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_167_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_167_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_167_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_167_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_167_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_167_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_167_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_167_8;
  wire                _zz_when_ArraySlice_l418_6;
  wire                _zz_when_ArraySlice_l418_6_1;
  wire                _zz_when_ArraySlice_l418_6_2;
  wire                _zz_when_ArraySlice_l418_6_3;
  wire                _zz_when_ArraySlice_l418_6_4;
  wire                _zz_when_ArraySlice_l418_6_5;
  wire       [5:0]    _zz_when_ArraySlice_l421_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l421_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l421_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l421_6_4;
  wire       [5:0]    _zz_when_ArraySlice_l421_6_5;
  wire       [0:0]    _zz_when_ArraySlice_l421_6_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_6_7;
  wire       [5:0]    _zz_selectReadFifo_6_24;
  wire       [0:0]    _zz_selectReadFifo_6_25;
  wire       [12:0]   _zz_when_ArraySlice_l425_6;
  wire       [12:0]   _zz_when_ArraySlice_l425_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l425_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l425_6_3;
  wire       [12:0]   _zz_when_ArraySlice_l436_6;
  wire       [5:0]    _zz_when_ArraySlice_l436_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l436_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l436_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l436_6_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_20;
  wire       [6:0]    _zz_when_ArraySlice_l95_20;
  wire       [6:0]    _zz_when_ArraySlice_l95_20_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_20_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_20_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_20_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_6;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_6_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_6_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_20;
  wire       [6:0]    _zz_when_ArraySlice_l99_20_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l437_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l437_6_4;
  wire       [5:0]    _zz_selectReadFifo_6_26;
  wire       [5:0]    _zz_selectReadFifo_6_27;
  wire       [5:0]    _zz_selectReadFifo_6_28;
  wire       [0:0]    _zz_selectReadFifo_6_29;
  wire       [5:0]    _zz_when_ArraySlice_l165_168;
  wire       [5:0]    _zz_when_ArraySlice_l165_168_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_168_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_168;
  wire       [6:0]    _zz_when_ArraySlice_l166_168_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_168_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_168_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_168_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_168_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_168;
  wire       [6:0]    _zz_when_ArraySlice_l113_168;
  wire       [6:0]    _zz_when_ArraySlice_l113_168_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_168_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_168_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_168_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_168;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_168_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_168_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_168_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_168;
  wire       [6:0]    _zz_when_ArraySlice_l118_168_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_168_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_168_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_168_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_168_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_168_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_168_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_168_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_168_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_169;
  wire       [5:0]    _zz_when_ArraySlice_l165_169_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_169_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_169;
  wire       [5:0]    _zz_when_ArraySlice_l166_169_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_169_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_169_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_169_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_169;
  wire       [6:0]    _zz_when_ArraySlice_l113_169;
  wire       [6:0]    _zz_when_ArraySlice_l113_169_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_169_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_169_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_169_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_169;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_169_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_169_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_169_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_169;
  wire       [6:0]    _zz_when_ArraySlice_l118_169_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_169_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_169_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_169_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_169_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_169_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_169_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_169_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_169_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_169_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_170;
  wire       [5:0]    _zz_when_ArraySlice_l165_170_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_170_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_170;
  wire       [5:0]    _zz_when_ArraySlice_l166_170_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_170_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_170_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_170_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_170;
  wire       [6:0]    _zz_when_ArraySlice_l113_170;
  wire       [6:0]    _zz_when_ArraySlice_l113_170_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_170_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_170_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_170_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_170;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_170_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_170_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_170_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_170;
  wire       [6:0]    _zz_when_ArraySlice_l118_170_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_170_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_170_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_170_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_170_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_170_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_170_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_170_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_170_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_170_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_171;
  wire       [5:0]    _zz_when_ArraySlice_l165_171_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_171_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_171;
  wire       [5:0]    _zz_when_ArraySlice_l166_171_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_171_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_171_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_171_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_171;
  wire       [6:0]    _zz_when_ArraySlice_l113_171;
  wire       [6:0]    _zz_when_ArraySlice_l113_171_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_171_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_171_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_171_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_171;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_171_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_171_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_171_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_171;
  wire       [6:0]    _zz_when_ArraySlice_l118_171_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_171_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_171_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_171_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_171_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_171_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_171_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_171_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_171_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_171_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_172;
  wire       [5:0]    _zz_when_ArraySlice_l165_172_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_172;
  wire       [5:0]    _zz_when_ArraySlice_l166_172_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_172_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_172_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_172;
  wire       [6:0]    _zz_when_ArraySlice_l113_172;
  wire       [6:0]    _zz_when_ArraySlice_l113_172_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_172_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_172_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_172_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_172;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_172_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_172_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_172_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_172;
  wire       [6:0]    _zz_when_ArraySlice_l118_172_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_172_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_172_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_172_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_172_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_172_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_172_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_172_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_172_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_173;
  wire       [5:0]    _zz_when_ArraySlice_l165_173_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_173;
  wire       [4:0]    _zz_when_ArraySlice_l166_173_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_173_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_173_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_173_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_173;
  wire       [6:0]    _zz_when_ArraySlice_l113_173;
  wire       [6:0]    _zz_when_ArraySlice_l113_173_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_173_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_173_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_173_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_173;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_173_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_173_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_173_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_173;
  wire       [6:0]    _zz_when_ArraySlice_l118_173_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_173_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_173_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_173_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_173_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_173_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_173_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_173_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_173_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_174;
  wire       [5:0]    _zz_when_ArraySlice_l165_174_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_174;
  wire       [4:0]    _zz_when_ArraySlice_l166_174_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_174_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_174_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_174_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_174;
  wire       [6:0]    _zz_when_ArraySlice_l113_174;
  wire       [6:0]    _zz_when_ArraySlice_l113_174_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_174_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_174_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_174_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_174;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_174_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_174_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_174_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_174;
  wire       [6:0]    _zz_when_ArraySlice_l118_174_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_174_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_174_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_174_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_174_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_174_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_174_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_174_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_174_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_175;
  wire       [5:0]    _zz_when_ArraySlice_l165_175_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_175;
  wire       [3:0]    _zz_when_ArraySlice_l166_175_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_175_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_175_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_175_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_175;
  wire       [6:0]    _zz_when_ArraySlice_l113_175;
  wire       [6:0]    _zz_when_ArraySlice_l113_175_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_175_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_175_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_175_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_175;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_175_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_175_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_175_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_175;
  wire       [6:0]    _zz_when_ArraySlice_l118_175_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_175_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_175_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_175_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_175_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_175_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_175_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_175_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_175_8;
  wire                _zz_when_ArraySlice_l444_6;
  wire                _zz_when_ArraySlice_l444_6_1;
  wire                _zz_when_ArraySlice_l444_6_2;
  wire                _zz_when_ArraySlice_l444_6_3;
  wire                _zz_when_ArraySlice_l444_6_4;
  wire                _zz_when_ArraySlice_l444_6_5;
  wire       [5:0]    _zz_selectReadFifo_6_30;
  wire       [0:0]    _zz_selectReadFifo_6_31;
  wire       [12:0]   _zz_when_ArraySlice_l448_6;
  wire       [12:0]   _zz_when_ArraySlice_l448_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l448_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l448_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l434_6;
  wire       [5:0]    _zz_when_ArraySlice_l434_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l455_6;
  wire       [5:0]    _zz_when_ArraySlice_l455_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l455_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l455_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l455_6_4;
  wire       [5:0]    _zz_when_ArraySlice_l373_7;
  wire       [5:0]    _zz_when_ArraySlice_l373_7_1;
  reg        [6:0]    _zz_when_ArraySlice_l374_7;
  wire       [5:0]    _zz_when_ArraySlice_l374_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l374_7_2;
  wire       [5:0]    _zz__zz_outputStreamArrayData_7_valid;
  reg                 _zz_outputStreamArrayData_7_valid_2;
  reg        [31:0]   _zz_outputStreamArrayData_7_payload;
  wire       [6:0]    _zz_when_ArraySlice_l380_7;
  wire       [0:0]    _zz_when_ArraySlice_l380_7_1;
  reg        [6:0]    _zz_when_ArraySlice_l380_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l380_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l380_7_4;
  wire       [12:0]   _zz_when_ArraySlice_l381_7;
  wire       [5:0]    _zz_when_ArraySlice_l381_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l381_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l381_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l381_7_4;
  wire       [5:0]    _zz_selectReadFifo_7;
  wire       [5:0]    _zz_selectReadFifo_7_1;
  wire       [5:0]    _zz_selectReadFifo_7_2;
  wire       [0:0]    _zz_selectReadFifo_7_3;
  wire       [5:0]    _zz_selectReadFifo_7_4;
  wire       [0:0]    _zz_selectReadFifo_7_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_7;
  wire       [12:0]   _zz_when_ArraySlice_l384_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l384_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l384_7_3;
  reg        [6:0]    _zz_when_ArraySlice_l389_7;
  wire       [5:0]    _zz_when_ArraySlice_l389_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l389_7_2;
  wire       [6:0]    _zz_when_ArraySlice_l389_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l389_7_4;
  wire       [12:0]   _zz_when_ArraySlice_l390_7;
  wire       [5:0]    _zz_when_ArraySlice_l390_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l390_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l390_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l390_7_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_21;
  wire       [6:0]    _zz_when_ArraySlice_l95_21;
  wire       [6:0]    _zz_when_ArraySlice_l95_21_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_21_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_21_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_21_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_7;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_7_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_7_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l392_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_21;
  wire       [6:0]    _zz_when_ArraySlice_l99_21_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l392_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l392_7_4;
  wire       [5:0]    _zz_selectReadFifo_7_6;
  wire       [5:0]    _zz_selectReadFifo_7_7;
  wire       [5:0]    _zz_selectReadFifo_7_8;
  wire       [0:0]    _zz_selectReadFifo_7_9;
  wire       [5:0]    _zz_selectReadFifo_7_10;
  wire       [5:0]    _zz_selectReadFifo_7_11;
  wire       [5:0]    _zz_selectReadFifo_7_12;
  wire       [0:0]    _zz_selectReadFifo_7_13;
  wire       [5:0]    _zz_when_ArraySlice_l165_176;
  wire       [5:0]    _zz_when_ArraySlice_l165_176_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_176_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_176;
  wire       [6:0]    _zz_when_ArraySlice_l166_176_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_176_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_176_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_176_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_176_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_176;
  wire       [6:0]    _zz_when_ArraySlice_l113_176;
  wire       [6:0]    _zz_when_ArraySlice_l113_176_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_176_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_176_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_176_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_176;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_176_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_176_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_176_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_176;
  wire       [6:0]    _zz_when_ArraySlice_l118_176_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_176_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_176_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_176_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_176_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_176_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_176_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_176_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_176_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_177;
  wire       [5:0]    _zz_when_ArraySlice_l165_177_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_177_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_177;
  wire       [5:0]    _zz_when_ArraySlice_l166_177_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_177_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_177_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_177_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_177;
  wire       [6:0]    _zz_when_ArraySlice_l113_177;
  wire       [6:0]    _zz_when_ArraySlice_l113_177_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_177_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_177_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_177_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_177;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_177_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_177_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_177_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_177;
  wire       [6:0]    _zz_when_ArraySlice_l118_177_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_177_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_177_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_177_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_177_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_177_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_177_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_177_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_177_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_177_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_178;
  wire       [5:0]    _zz_when_ArraySlice_l165_178_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_178_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_178;
  wire       [5:0]    _zz_when_ArraySlice_l166_178_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_178_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_178_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_178_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_178;
  wire       [6:0]    _zz_when_ArraySlice_l113_178;
  wire       [6:0]    _zz_when_ArraySlice_l113_178_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_178_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_178_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_178_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_178;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_178_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_178_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_178_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_178;
  wire       [6:0]    _zz_when_ArraySlice_l118_178_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_178_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_178_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_178_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_178_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_178_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_178_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_178_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_178_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_178_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_179;
  wire       [5:0]    _zz_when_ArraySlice_l165_179_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_179_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_179;
  wire       [5:0]    _zz_when_ArraySlice_l166_179_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_179_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_179_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_179_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_179;
  wire       [6:0]    _zz_when_ArraySlice_l113_179;
  wire       [6:0]    _zz_when_ArraySlice_l113_179_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_179_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_179_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_179_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_179;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_179_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_179_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_179_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_179;
  wire       [6:0]    _zz_when_ArraySlice_l118_179_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_179_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_179_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_179_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_179_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_179_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_179_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_179_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_179_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_179_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_180;
  wire       [5:0]    _zz_when_ArraySlice_l165_180_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_180;
  wire       [5:0]    _zz_when_ArraySlice_l166_180_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_180_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_180_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_180;
  wire       [6:0]    _zz_when_ArraySlice_l113_180;
  wire       [6:0]    _zz_when_ArraySlice_l113_180_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_180_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_180_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_180_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_180;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_180_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_180_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_180_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_180;
  wire       [6:0]    _zz_when_ArraySlice_l118_180_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_180_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_180_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_180_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_180_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_180_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_180_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_180_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_180_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_181;
  wire       [5:0]    _zz_when_ArraySlice_l165_181_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_181;
  wire       [4:0]    _zz_when_ArraySlice_l166_181_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_181_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_181_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_181_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_181;
  wire       [6:0]    _zz_when_ArraySlice_l113_181;
  wire       [6:0]    _zz_when_ArraySlice_l113_181_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_181_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_181_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_181_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_181;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_181_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_181_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_181_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_181;
  wire       [6:0]    _zz_when_ArraySlice_l118_181_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_181_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_181_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_181_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_181_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_181_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_181_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_181_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_181_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_182;
  wire       [5:0]    _zz_when_ArraySlice_l165_182_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_182;
  wire       [4:0]    _zz_when_ArraySlice_l166_182_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_182_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_182_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_182_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_182;
  wire       [6:0]    _zz_when_ArraySlice_l113_182;
  wire       [6:0]    _zz_when_ArraySlice_l113_182_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_182_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_182_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_182_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_182;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_182_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_182_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_182_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_182;
  wire       [6:0]    _zz_when_ArraySlice_l118_182_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_182_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_182_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_182_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_182_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_182_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_182_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_182_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_182_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_183;
  wire       [5:0]    _zz_when_ArraySlice_l165_183_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_183;
  wire       [3:0]    _zz_when_ArraySlice_l166_183_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_183_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_183_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_183_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_183;
  wire       [6:0]    _zz_when_ArraySlice_l113_183;
  wire       [6:0]    _zz_when_ArraySlice_l113_183_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_183_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_183_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_183_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_183;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_183_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_183_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_183_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_183;
  wire       [6:0]    _zz_when_ArraySlice_l118_183_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_183_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_183_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_183_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_183_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_183_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_183_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_183_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_183_8;
  wire                _zz_when_ArraySlice_l398_7_1;
  wire                _zz_when_ArraySlice_l398_7_2;
  wire                _zz_when_ArraySlice_l398_7_3;
  wire                _zz_when_ArraySlice_l398_7_4;
  wire                _zz_when_ArraySlice_l398_7_5;
  wire                _zz_when_ArraySlice_l398_7_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l401_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l401_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l401_7_4;
  wire       [5:0]    _zz_when_ArraySlice_l401_7_5;
  wire       [0:0]    _zz_when_ArraySlice_l401_7_6;
  wire       [5:0]    _zz_when_ArraySlice_l401_7_7;
  wire       [5:0]    _zz_selectReadFifo_7_14;
  wire       [0:0]    _zz_selectReadFifo_7_15;
  wire       [12:0]   _zz_when_ArraySlice_l405_7;
  wire       [12:0]   _zz_when_ArraySlice_l405_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l405_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l405_7_3;
  reg        [6:0]    _zz_when_ArraySlice_l409_7;
  wire       [5:0]    _zz_when_ArraySlice_l409_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l409_7_2;
  wire       [12:0]   _zz_when_ArraySlice_l410_7;
  wire       [5:0]    _zz_when_ArraySlice_l410_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l410_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l410_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l410_7_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_22;
  wire       [6:0]    _zz_when_ArraySlice_l95_22;
  wire       [6:0]    _zz_when_ArraySlice_l95_22_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_22_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_22_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_22_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_7;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_7_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_7_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l412_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_22;
  wire       [6:0]    _zz_when_ArraySlice_l99_22_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l412_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l412_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l412_7_4;
  wire       [5:0]    _zz_selectReadFifo_7_16;
  wire       [5:0]    _zz_selectReadFifo_7_17;
  wire       [5:0]    _zz_selectReadFifo_7_18;
  wire       [0:0]    _zz_selectReadFifo_7_19;
  wire       [5:0]    _zz_selectReadFifo_7_20;
  wire       [5:0]    _zz_selectReadFifo_7_21;
  wire       [5:0]    _zz_selectReadFifo_7_22;
  wire       [0:0]    _zz_selectReadFifo_7_23;
  wire       [5:0]    _zz_when_ArraySlice_l165_184;
  wire       [5:0]    _zz_when_ArraySlice_l165_184_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_184_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_184;
  wire       [6:0]    _zz_when_ArraySlice_l166_184_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_184_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_184_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_184_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_184_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_184;
  wire       [6:0]    _zz_when_ArraySlice_l113_184;
  wire       [6:0]    _zz_when_ArraySlice_l113_184_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_184_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_184_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_184_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_184;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_184_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_184_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_184_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_184;
  wire       [6:0]    _zz_when_ArraySlice_l118_184_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_184_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_184_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_184_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_184_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_184_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_184_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_184_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_184_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_185;
  wire       [5:0]    _zz_when_ArraySlice_l165_185_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_185_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_185;
  wire       [5:0]    _zz_when_ArraySlice_l166_185_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_185_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_185_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_185_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_185;
  wire       [6:0]    _zz_when_ArraySlice_l113_185;
  wire       [6:0]    _zz_when_ArraySlice_l113_185_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_185_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_185_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_185_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_185;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_185_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_185_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_185_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_185;
  wire       [6:0]    _zz_when_ArraySlice_l118_185_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_185_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_185_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_185_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_185_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_185_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_185_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_185_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_185_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_185_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_186;
  wire       [5:0]    _zz_when_ArraySlice_l165_186_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_186_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_186;
  wire       [5:0]    _zz_when_ArraySlice_l166_186_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_186_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_186_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_186_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_186;
  wire       [6:0]    _zz_when_ArraySlice_l113_186;
  wire       [6:0]    _zz_when_ArraySlice_l113_186_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_186_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_186_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_186_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_186;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_186_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_186_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_186_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_186;
  wire       [6:0]    _zz_when_ArraySlice_l118_186_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_186_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_186_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_186_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_186_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_186_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_186_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_186_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_186_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_186_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_187;
  wire       [5:0]    _zz_when_ArraySlice_l165_187_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_187_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_187;
  wire       [5:0]    _zz_when_ArraySlice_l166_187_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_187_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_187_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_187_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_187;
  wire       [6:0]    _zz_when_ArraySlice_l113_187;
  wire       [6:0]    _zz_when_ArraySlice_l113_187_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_187_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_187_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_187_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_187;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_187_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_187_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_187_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_187;
  wire       [6:0]    _zz_when_ArraySlice_l118_187_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_187_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_187_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_187_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_187_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_187_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_187_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_187_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_187_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_187_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_188;
  wire       [5:0]    _zz_when_ArraySlice_l165_188_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_188;
  wire       [5:0]    _zz_when_ArraySlice_l166_188_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_188_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_188_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_188;
  wire       [6:0]    _zz_when_ArraySlice_l113_188;
  wire       [6:0]    _zz_when_ArraySlice_l113_188_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_188_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_188_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_188_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_188;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_188_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_188_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_188_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_188;
  wire       [6:0]    _zz_when_ArraySlice_l118_188_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_188_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_188_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_188_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_188_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_188_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_188_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_188_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_188_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_189;
  wire       [5:0]    _zz_when_ArraySlice_l165_189_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_189;
  wire       [4:0]    _zz_when_ArraySlice_l166_189_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_189_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_189_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_189_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_189;
  wire       [6:0]    _zz_when_ArraySlice_l113_189;
  wire       [6:0]    _zz_when_ArraySlice_l113_189_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_189_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_189_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_189_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_189;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_189_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_189_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_189_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_189;
  wire       [6:0]    _zz_when_ArraySlice_l118_189_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_189_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_189_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_189_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_189_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_189_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_189_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_189_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_189_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_190;
  wire       [5:0]    _zz_when_ArraySlice_l165_190_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_190;
  wire       [4:0]    _zz_when_ArraySlice_l166_190_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_190_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_190_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_190_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_190;
  wire       [6:0]    _zz_when_ArraySlice_l113_190;
  wire       [6:0]    _zz_when_ArraySlice_l113_190_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_190_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_190_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_190_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_190;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_190_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_190_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_190_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_190;
  wire       [6:0]    _zz_when_ArraySlice_l118_190_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_190_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_190_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_190_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_190_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_190_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_190_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_190_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_190_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_191;
  wire       [5:0]    _zz_when_ArraySlice_l165_191_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_191;
  wire       [3:0]    _zz_when_ArraySlice_l166_191_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_191_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_191_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_191_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_191;
  wire       [6:0]    _zz_when_ArraySlice_l113_191;
  wire       [6:0]    _zz_when_ArraySlice_l113_191_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_191_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_191_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_191_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_191;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_191_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_191_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_191_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_191;
  wire       [6:0]    _zz_when_ArraySlice_l118_191_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_191_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_191_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_191_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_191_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_191_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_191_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_191_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_191_8;
  wire                _zz_when_ArraySlice_l418_7;
  wire                _zz_when_ArraySlice_l418_7_1;
  wire                _zz_when_ArraySlice_l418_7_2;
  wire                _zz_when_ArraySlice_l418_7_3;
  wire                _zz_when_ArraySlice_l418_7_4;
  wire                _zz_when_ArraySlice_l418_7_5;
  wire       [5:0]    _zz_when_ArraySlice_l421_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l421_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l421_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l421_7_4;
  wire       [5:0]    _zz_when_ArraySlice_l421_7_5;
  wire       [0:0]    _zz_when_ArraySlice_l421_7_6;
  wire       [5:0]    _zz_when_ArraySlice_l421_7_7;
  wire       [5:0]    _zz_selectReadFifo_7_24;
  wire       [0:0]    _zz_selectReadFifo_7_25;
  wire       [12:0]   _zz_when_ArraySlice_l425_7;
  wire       [12:0]   _zz_when_ArraySlice_l425_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l425_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l425_7_3;
  wire       [12:0]   _zz_when_ArraySlice_l436_7;
  wire       [5:0]    _zz_when_ArraySlice_l436_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l436_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l436_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l436_7_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_23;
  wire       [6:0]    _zz_when_ArraySlice_l95_23;
  wire       [6:0]    _zz_when_ArraySlice_l95_23_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_23_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_23_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_23_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_7;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_7_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_7_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l437_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_23;
  wire       [6:0]    _zz_when_ArraySlice_l99_23_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l437_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l437_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l437_7_4;
  wire       [5:0]    _zz_selectReadFifo_7_26;
  wire       [5:0]    _zz_selectReadFifo_7_27;
  wire       [5:0]    _zz_selectReadFifo_7_28;
  wire       [0:0]    _zz_selectReadFifo_7_29;
  wire       [5:0]    _zz_when_ArraySlice_l165_192;
  wire       [5:0]    _zz_when_ArraySlice_l165_192_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_192_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_192;
  wire       [6:0]    _zz_when_ArraySlice_l166_192_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_192_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_192_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_192_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_192_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_192;
  wire       [6:0]    _zz_when_ArraySlice_l113_192;
  wire       [6:0]    _zz_when_ArraySlice_l113_192_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_192_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_192_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_192_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_192;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_192_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_192_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_192_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_192;
  wire       [6:0]    _zz_when_ArraySlice_l118_192_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_192_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_192_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_192_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_192_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_192_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_192_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_192_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_192_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_193;
  wire       [5:0]    _zz_when_ArraySlice_l165_193_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_193_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_193;
  wire       [5:0]    _zz_when_ArraySlice_l166_193_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_193_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_193_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_193_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_193;
  wire       [6:0]    _zz_when_ArraySlice_l113_193;
  wire       [6:0]    _zz_when_ArraySlice_l113_193_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_193_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_193_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_193_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_193;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_193_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_193_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_193_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_193;
  wire       [6:0]    _zz_when_ArraySlice_l118_193_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_193_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_193_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_193_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_193_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_193_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_193_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_193_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_193_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_193_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_194;
  wire       [5:0]    _zz_when_ArraySlice_l165_194_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_194_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_194;
  wire       [5:0]    _zz_when_ArraySlice_l166_194_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_194_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_194_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_194_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_194;
  wire       [6:0]    _zz_when_ArraySlice_l113_194;
  wire       [6:0]    _zz_when_ArraySlice_l113_194_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_194_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_194_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_194_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_194;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_194_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_194_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_194_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_194;
  wire       [6:0]    _zz_when_ArraySlice_l118_194_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_194_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_194_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_194_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_194_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_194_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_194_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_194_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_194_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_194_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_195;
  wire       [5:0]    _zz_when_ArraySlice_l165_195_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_195_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_195;
  wire       [5:0]    _zz_when_ArraySlice_l166_195_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_195_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_195_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_195_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_195;
  wire       [6:0]    _zz_when_ArraySlice_l113_195;
  wire       [6:0]    _zz_when_ArraySlice_l113_195_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_195_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_195_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_195_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_195;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_195_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_195_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_195_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_195;
  wire       [6:0]    _zz_when_ArraySlice_l118_195_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_195_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_195_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_195_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_195_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_195_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_195_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_195_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_195_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_195_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_196;
  wire       [5:0]    _zz_when_ArraySlice_l165_196_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_196;
  wire       [5:0]    _zz_when_ArraySlice_l166_196_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_196_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_196_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_196;
  wire       [6:0]    _zz_when_ArraySlice_l113_196;
  wire       [6:0]    _zz_when_ArraySlice_l113_196_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_196_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_196_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_196_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_196;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_196_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_196_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_196_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_196;
  wire       [6:0]    _zz_when_ArraySlice_l118_196_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_196_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_196_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_196_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_196_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_196_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_196_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_196_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_196_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_197;
  wire       [5:0]    _zz_when_ArraySlice_l165_197_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_197;
  wire       [4:0]    _zz_when_ArraySlice_l166_197_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_197_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_197_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_197_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_197;
  wire       [6:0]    _zz_when_ArraySlice_l113_197;
  wire       [6:0]    _zz_when_ArraySlice_l113_197_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_197_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_197_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_197_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_197;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_197_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_197_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_197_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_197;
  wire       [6:0]    _zz_when_ArraySlice_l118_197_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_197_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_197_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_197_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_197_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_197_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_197_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_197_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_197_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_198;
  wire       [5:0]    _zz_when_ArraySlice_l165_198_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_198;
  wire       [4:0]    _zz_when_ArraySlice_l166_198_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_198_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_198_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_198_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_198;
  wire       [6:0]    _zz_when_ArraySlice_l113_198;
  wire       [6:0]    _zz_when_ArraySlice_l113_198_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_198_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_198_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_198_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_198;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_198_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_198_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_198_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_198;
  wire       [6:0]    _zz_when_ArraySlice_l118_198_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_198_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_198_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_198_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_198_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_198_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_198_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_198_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_198_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_199;
  wire       [5:0]    _zz_when_ArraySlice_l165_199_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_199;
  wire       [3:0]    _zz_when_ArraySlice_l166_199_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_199_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_199_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_199_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_199;
  wire       [6:0]    _zz_when_ArraySlice_l113_199;
  wire       [6:0]    _zz_when_ArraySlice_l113_199_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_199_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_199_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_199_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_199;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_199_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_199_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_199_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_199;
  wire       [6:0]    _zz_when_ArraySlice_l118_199_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_199_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_199_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_199_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_199_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_199_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_199_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_199_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_199_8;
  wire                _zz_when_ArraySlice_l444_7;
  wire                _zz_when_ArraySlice_l444_7_1;
  wire                _zz_when_ArraySlice_l444_7_2;
  wire                _zz_when_ArraySlice_l444_7_3;
  wire                _zz_when_ArraySlice_l444_7_4;
  wire                _zz_when_ArraySlice_l444_7_5;
  wire       [5:0]    _zz_selectReadFifo_7_30;
  wire       [0:0]    _zz_selectReadFifo_7_31;
  wire       [12:0]   _zz_when_ArraySlice_l448_7;
  wire       [12:0]   _zz_when_ArraySlice_l448_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l448_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l448_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l434_7;
  wire       [5:0]    _zz_when_ArraySlice_l434_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l455_7;
  wire       [5:0]    _zz_when_ArraySlice_l455_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l455_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l455_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l455_7_4;
  wire       [5:0]    _zz_when_ArraySlice_l165_200;
  wire       [5:0]    _zz_when_ArraySlice_l165_200_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_200_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_200;
  wire       [6:0]    _zz_when_ArraySlice_l166_200_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_200_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_200_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_200_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_200_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_200;
  wire       [6:0]    _zz_when_ArraySlice_l113_200;
  wire       [6:0]    _zz_when_ArraySlice_l113_200_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_200_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_200_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_200_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_200;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_200_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_200_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_200_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_200;
  wire       [6:0]    _zz_when_ArraySlice_l118_200_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_200_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_200_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_200_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_200_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_200_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_200_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_200_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_200_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_201;
  wire       [5:0]    _zz_when_ArraySlice_l165_201_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_201_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_201;
  wire       [5:0]    _zz_when_ArraySlice_l166_201_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_201_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_201_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_201_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_201;
  wire       [6:0]    _zz_when_ArraySlice_l113_201;
  wire       [6:0]    _zz_when_ArraySlice_l113_201_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_201_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_201_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_201_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_201;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_201_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_201_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_201_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_201;
  wire       [6:0]    _zz_when_ArraySlice_l118_201_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_201_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_201_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_201_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_201_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_201_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_201_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_201_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_201_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_201_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_202;
  wire       [5:0]    _zz_when_ArraySlice_l165_202_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_202_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_202;
  wire       [5:0]    _zz_when_ArraySlice_l166_202_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_202_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_202_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_202_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_202;
  wire       [6:0]    _zz_when_ArraySlice_l113_202;
  wire       [6:0]    _zz_when_ArraySlice_l113_202_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_202_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_202_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_202_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_202;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_202_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_202_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_202_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_202;
  wire       [6:0]    _zz_when_ArraySlice_l118_202_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_202_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_202_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_202_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_202_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_202_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_202_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_202_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_202_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_202_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_203;
  wire       [5:0]    _zz_when_ArraySlice_l165_203_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_203_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_203;
  wire       [5:0]    _zz_when_ArraySlice_l166_203_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_203_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_203_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_203_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_203;
  wire       [6:0]    _zz_when_ArraySlice_l113_203;
  wire       [6:0]    _zz_when_ArraySlice_l113_203_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_203_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_203_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_203_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_203;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_203_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_203_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_203_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_203;
  wire       [6:0]    _zz_when_ArraySlice_l118_203_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_203_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_203_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_203_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_203_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_203_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_203_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_203_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_203_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_203_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_204;
  wire       [5:0]    _zz_when_ArraySlice_l165_204_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_204;
  wire       [5:0]    _zz_when_ArraySlice_l166_204_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_204_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_204_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_204;
  wire       [6:0]    _zz_when_ArraySlice_l113_204;
  wire       [6:0]    _zz_when_ArraySlice_l113_204_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_204_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_204_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_204_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_204;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_204_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_204_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_204_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_204;
  wire       [6:0]    _zz_when_ArraySlice_l118_204_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_204_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_204_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_204_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_204_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_204_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_204_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_204_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_204_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_205;
  wire       [5:0]    _zz_when_ArraySlice_l165_205_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_205;
  wire       [4:0]    _zz_when_ArraySlice_l166_205_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_205_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_205_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_205_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_205;
  wire       [6:0]    _zz_when_ArraySlice_l113_205;
  wire       [6:0]    _zz_when_ArraySlice_l113_205_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_205_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_205_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_205_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_205;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_205_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_205_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_205_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_205;
  wire       [6:0]    _zz_when_ArraySlice_l118_205_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_205_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_205_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_205_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_205_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_205_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_205_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_205_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_205_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_206;
  wire       [5:0]    _zz_when_ArraySlice_l165_206_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_206;
  wire       [4:0]    _zz_when_ArraySlice_l166_206_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_206_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_206_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_206_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_206;
  wire       [6:0]    _zz_when_ArraySlice_l113_206;
  wire       [6:0]    _zz_when_ArraySlice_l113_206_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_206_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_206_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_206_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_206;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_206_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_206_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_206_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_206;
  wire       [6:0]    _zz_when_ArraySlice_l118_206_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_206_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_206_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_206_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_206_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_206_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_206_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_206_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_206_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_207;
  wire       [5:0]    _zz_when_ArraySlice_l165_207_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_207;
  wire       [3:0]    _zz_when_ArraySlice_l166_207_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_207_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_207_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_207_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_207;
  wire       [6:0]    _zz_when_ArraySlice_l113_207;
  wire       [6:0]    _zz_when_ArraySlice_l113_207_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_207_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_207_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_207_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_207;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_207_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_207_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_207_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_207;
  wire       [6:0]    _zz_when_ArraySlice_l118_207_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_207_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_207_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_207_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_207_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_207_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_207_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_207_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_207_8;
  wire                _zz_when_ArraySlice_l465;
  wire                _zz_when_ArraySlice_l465_1;
  wire                _zz_when_ArraySlice_l465_2;
  wire                _zz_when_ArraySlice_l465_3;
  wire                _zz_when_ArraySlice_l465_4;
  wire                _zz_when_ArraySlice_l465_5;
  wire       [5:0]    _zz_when_ArraySlice_l240;
  wire       [5:0]    _zz_when_ArraySlice_l240_1;
  wire       [2:0]    _zz_when_ArraySlice_l240_2;
  reg        [6:0]    _zz_when_ArraySlice_l241;
  wire       [5:0]    _zz_when_ArraySlice_l241_1;
  wire       [5:0]    _zz_when_ArraySlice_l241_2;
  wire       [2:0]    _zz_when_ArraySlice_l241_3;
  wire       [5:0]    _zz__zz_outputStreamArrayData_0_valid_1_1;
  wire       [2:0]    _zz__zz_outputStreamArrayData_0_valid_1_2;
  reg                 _zz_outputStreamArrayData_0_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_0_payload_1;
  wire       [6:0]    _zz_when_ArraySlice_l247;
  wire       [0:0]    _zz_when_ArraySlice_l247_1;
  reg        [6:0]    _zz_when_ArraySlice_l247_2;
  wire       [5:0]    _zz_when_ArraySlice_l247_3;
  wire       [5:0]    _zz_when_ArraySlice_l247_4;
  wire       [2:0]    _zz_when_ArraySlice_l247_5;
  wire       [12:0]   _zz_when_ArraySlice_l248;
  wire       [5:0]    _zz_when_ArraySlice_l248_1;
  wire       [5:0]    _zz_when_ArraySlice_l248_2;
  wire       [5:0]    _zz_when_ArraySlice_l248_3;
  wire       [0:0]    _zz_when_ArraySlice_l248_4;
  wire       [5:0]    _zz_selectReadFifo_0_32;
  wire       [5:0]    _zz_selectReadFifo_0_33;
  wire       [5:0]    _zz_selectReadFifo_0_34;
  wire       [0:0]    _zz_selectReadFifo_0_35;
  wire       [5:0]    _zz_selectReadFifo_0_36;
  wire       [0:0]    _zz_selectReadFifo_0_37;
  wire       [12:0]   _zz_when_ArraySlice_l251;
  wire       [12:0]   _zz_when_ArraySlice_l251_1;
  wire       [12:0]   _zz_when_ArraySlice_l251_2;
  wire       [0:0]    _zz_when_ArraySlice_l251_3;
  reg        [6:0]    _zz_when_ArraySlice_l256;
  wire       [5:0]    _zz_when_ArraySlice_l256_1;
  wire       [5:0]    _zz_when_ArraySlice_l256_2;
  wire       [2:0]    _zz_when_ArraySlice_l256_3;
  wire       [6:0]    _zz_when_ArraySlice_l256_4;
  wire       [0:0]    _zz_when_ArraySlice_l256_5;
  wire       [12:0]   _zz_when_ArraySlice_l257;
  wire       [5:0]    _zz_when_ArraySlice_l257_1;
  wire       [5:0]    _zz_when_ArraySlice_l257_2;
  wire       [5:0]    _zz_when_ArraySlice_l257_3;
  wire       [0:0]    _zz_when_ArraySlice_l257_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_24;
  wire       [6:0]    _zz_when_ArraySlice_l95_24;
  wire       [6:0]    _zz_when_ArraySlice_l95_24_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_24_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_24_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_24_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_24;
  wire       [6:0]    _zz_when_ArraySlice_l99_24_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_8;
  wire       [6:0]    _zz_when_ArraySlice_l259_9;
  wire       [0:0]    _zz_when_ArraySlice_l259_10;
  wire       [6:0]    _zz_when_ArraySlice_l259_11;
  wire       [5:0]    _zz_selectReadFifo_0_38;
  wire       [5:0]    _zz_selectReadFifo_0_39;
  wire       [5:0]    _zz_selectReadFifo_0_40;
  wire       [0:0]    _zz_selectReadFifo_0_41;
  wire       [5:0]    _zz_selectReadFifo_0_42;
  wire       [5:0]    _zz_selectReadFifo_0_43;
  wire       [5:0]    _zz_selectReadFifo_0_44;
  wire       [0:0]    _zz_selectReadFifo_0_45;
  wire       [5:0]    _zz_when_ArraySlice_l165_208;
  wire       [5:0]    _zz_when_ArraySlice_l165_208_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_208_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_208;
  wire       [6:0]    _zz_when_ArraySlice_l166_208_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_208_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_208_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_208_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_208_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_208;
  wire       [6:0]    _zz_when_ArraySlice_l113_208;
  wire       [6:0]    _zz_when_ArraySlice_l113_208_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_208_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_208_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_208_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_208;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_208_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_208_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_208_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_208;
  wire       [6:0]    _zz_when_ArraySlice_l118_208_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_208_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_208_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_208_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_208_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_208_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_208_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_208_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_208_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_209;
  wire       [5:0]    _zz_when_ArraySlice_l165_209_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_209_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_209;
  wire       [5:0]    _zz_when_ArraySlice_l166_209_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_209_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_209_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_209_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_209;
  wire       [6:0]    _zz_when_ArraySlice_l113_209;
  wire       [6:0]    _zz_when_ArraySlice_l113_209_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_209_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_209_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_209_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_209;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_209_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_209_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_209_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_209;
  wire       [6:0]    _zz_when_ArraySlice_l118_209_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_209_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_209_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_209_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_209_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_209_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_209_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_209_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_209_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_209_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_210;
  wire       [5:0]    _zz_when_ArraySlice_l165_210_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_210_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_210;
  wire       [5:0]    _zz_when_ArraySlice_l166_210_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_210_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_210_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_210_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_210;
  wire       [6:0]    _zz_when_ArraySlice_l113_210;
  wire       [6:0]    _zz_when_ArraySlice_l113_210_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_210_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_210_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_210_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_210;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_210_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_210_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_210_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_210;
  wire       [6:0]    _zz_when_ArraySlice_l118_210_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_210_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_210_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_210_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_210_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_210_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_210_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_210_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_210_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_210_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_211;
  wire       [5:0]    _zz_when_ArraySlice_l165_211_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_211_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_211;
  wire       [5:0]    _zz_when_ArraySlice_l166_211_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_211_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_211_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_211_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_211;
  wire       [6:0]    _zz_when_ArraySlice_l113_211;
  wire       [6:0]    _zz_when_ArraySlice_l113_211_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_211_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_211_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_211_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_211;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_211_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_211_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_211_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_211;
  wire       [6:0]    _zz_when_ArraySlice_l118_211_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_211_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_211_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_211_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_211_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_211_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_211_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_211_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_211_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_211_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_212;
  wire       [5:0]    _zz_when_ArraySlice_l165_212_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_212;
  wire       [5:0]    _zz_when_ArraySlice_l166_212_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_212_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_212_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_212;
  wire       [6:0]    _zz_when_ArraySlice_l113_212;
  wire       [6:0]    _zz_when_ArraySlice_l113_212_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_212_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_212_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_212_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_212;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_212_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_212_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_212_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_212;
  wire       [6:0]    _zz_when_ArraySlice_l118_212_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_212_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_212_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_212_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_212_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_212_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_212_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_212_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_212_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_213;
  wire       [5:0]    _zz_when_ArraySlice_l165_213_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_213;
  wire       [4:0]    _zz_when_ArraySlice_l166_213_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_213_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_213_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_213_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_213;
  wire       [6:0]    _zz_when_ArraySlice_l113_213;
  wire       [6:0]    _zz_when_ArraySlice_l113_213_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_213_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_213_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_213_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_213;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_213_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_213_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_213_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_213;
  wire       [6:0]    _zz_when_ArraySlice_l118_213_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_213_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_213_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_213_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_213_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_213_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_213_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_213_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_213_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_214;
  wire       [5:0]    _zz_when_ArraySlice_l165_214_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_214;
  wire       [4:0]    _zz_when_ArraySlice_l166_214_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_214_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_214_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_214_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_214;
  wire       [6:0]    _zz_when_ArraySlice_l113_214;
  wire       [6:0]    _zz_when_ArraySlice_l113_214_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_214_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_214_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_214_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_214;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_214_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_214_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_214_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_214;
  wire       [6:0]    _zz_when_ArraySlice_l118_214_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_214_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_214_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_214_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_214_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_214_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_214_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_214_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_214_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_215;
  wire       [5:0]    _zz_when_ArraySlice_l165_215_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_215;
  wire       [3:0]    _zz_when_ArraySlice_l166_215_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_215_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_215_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_215_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_215;
  wire       [6:0]    _zz_when_ArraySlice_l113_215;
  wire       [6:0]    _zz_when_ArraySlice_l113_215_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_215_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_215_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_215_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_215;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_215_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_215_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_215_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_215;
  wire       [6:0]    _zz_when_ArraySlice_l118_215_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_215_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_215_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_215_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_215_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_215_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_215_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_215_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_215_8;
  wire                _zz_when_ArraySlice_l265;
  wire                _zz_when_ArraySlice_l265_1;
  wire                _zz_when_ArraySlice_l265_2;
  wire                _zz_when_ArraySlice_l265_3;
  wire                _zz_when_ArraySlice_l265_4;
  wire                _zz_when_ArraySlice_l265_5;
  wire       [5:0]    _zz_when_ArraySlice_l268;
  wire       [5:0]    _zz_when_ArraySlice_l268_1;
  wire       [5:0]    _zz_when_ArraySlice_l268_2;
  wire       [5:0]    _zz_when_ArraySlice_l268_3;
  wire       [5:0]    _zz_when_ArraySlice_l268_4;
  wire       [0:0]    _zz_when_ArraySlice_l268_5;
  wire       [5:0]    _zz_when_ArraySlice_l268_6;
  wire       [2:0]    _zz_when_ArraySlice_l268_7;
  wire       [5:0]    _zz_selectReadFifo_0_46;
  wire       [0:0]    _zz_selectReadFifo_0_47;
  wire       [12:0]   _zz_when_ArraySlice_l272;
  wire       [12:0]   _zz_when_ArraySlice_l272_1;
  wire       [12:0]   _zz_when_ArraySlice_l272_2;
  wire       [0:0]    _zz_when_ArraySlice_l272_3;
  reg        [6:0]    _zz_when_ArraySlice_l276;
  wire       [5:0]    _zz_when_ArraySlice_l276_1;
  wire       [5:0]    _zz_when_ArraySlice_l276_2;
  wire       [2:0]    _zz_when_ArraySlice_l276_3;
  wire       [12:0]   _zz_when_ArraySlice_l277;
  wire       [5:0]    _zz_when_ArraySlice_l277_1;
  wire       [5:0]    _zz_when_ArraySlice_l277_2;
  wire       [5:0]    _zz_when_ArraySlice_l277_3;
  wire       [0:0]    _zz_when_ArraySlice_l277_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_25;
  wire       [6:0]    _zz_when_ArraySlice_l95_25;
  wire       [6:0]    _zz_when_ArraySlice_l95_25_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_25_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_25_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_25_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_25;
  wire       [6:0]    _zz_when_ArraySlice_l99_25_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_8;
  wire       [6:0]    _zz_when_ArraySlice_l279_9;
  wire       [0:0]    _zz_when_ArraySlice_l279_10;
  wire       [6:0]    _zz_when_ArraySlice_l279_11;
  wire       [5:0]    _zz_selectReadFifo_0_48;
  wire       [5:0]    _zz_selectReadFifo_0_49;
  wire       [5:0]    _zz_selectReadFifo_0_50;
  wire       [0:0]    _zz_selectReadFifo_0_51;
  wire       [5:0]    _zz_selectReadFifo_0_52;
  wire       [5:0]    _zz_selectReadFifo_0_53;
  wire       [5:0]    _zz_selectReadFifo_0_54;
  wire       [0:0]    _zz_selectReadFifo_0_55;
  wire       [5:0]    _zz_when_ArraySlice_l165_216;
  wire       [5:0]    _zz_when_ArraySlice_l165_216_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_216_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_216;
  wire       [6:0]    _zz_when_ArraySlice_l166_216_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_216_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_216_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_216_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_216_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_216;
  wire       [6:0]    _zz_when_ArraySlice_l113_216;
  wire       [6:0]    _zz_when_ArraySlice_l113_216_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_216_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_216_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_216_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_216;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_216_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_216_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_216_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_216;
  wire       [6:0]    _zz_when_ArraySlice_l118_216_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_216_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_216_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_216_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_216_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_216_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_216_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_216_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_216_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_217;
  wire       [5:0]    _zz_when_ArraySlice_l165_217_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_217_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_217;
  wire       [5:0]    _zz_when_ArraySlice_l166_217_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_217_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_217_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_217_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_217;
  wire       [6:0]    _zz_when_ArraySlice_l113_217;
  wire       [6:0]    _zz_when_ArraySlice_l113_217_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_217_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_217_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_217_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_217;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_217_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_217_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_217_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_217;
  wire       [6:0]    _zz_when_ArraySlice_l118_217_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_217_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_217_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_217_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_217_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_217_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_217_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_217_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_217_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_217_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_218;
  wire       [5:0]    _zz_when_ArraySlice_l165_218_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_218_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_218;
  wire       [5:0]    _zz_when_ArraySlice_l166_218_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_218_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_218_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_218_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_218;
  wire       [6:0]    _zz_when_ArraySlice_l113_218;
  wire       [6:0]    _zz_when_ArraySlice_l113_218_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_218_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_218_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_218_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_218;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_218_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_218_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_218_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_218;
  wire       [6:0]    _zz_when_ArraySlice_l118_218_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_218_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_218_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_218_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_218_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_218_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_218_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_218_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_218_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_218_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_219;
  wire       [5:0]    _zz_when_ArraySlice_l165_219_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_219_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_219;
  wire       [5:0]    _zz_when_ArraySlice_l166_219_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_219_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_219_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_219_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_219;
  wire       [6:0]    _zz_when_ArraySlice_l113_219;
  wire       [6:0]    _zz_when_ArraySlice_l113_219_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_219_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_219_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_219_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_219;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_219_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_219_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_219_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_219;
  wire       [6:0]    _zz_when_ArraySlice_l118_219_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_219_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_219_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_219_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_219_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_219_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_219_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_219_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_219_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_219_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_220;
  wire       [5:0]    _zz_when_ArraySlice_l165_220_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_220;
  wire       [5:0]    _zz_when_ArraySlice_l166_220_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_220_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_220_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_220;
  wire       [6:0]    _zz_when_ArraySlice_l113_220;
  wire       [6:0]    _zz_when_ArraySlice_l113_220_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_220_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_220_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_220_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_220;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_220_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_220_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_220_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_220;
  wire       [6:0]    _zz_when_ArraySlice_l118_220_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_220_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_220_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_220_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_220_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_220_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_220_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_220_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_220_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_221;
  wire       [5:0]    _zz_when_ArraySlice_l165_221_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_221;
  wire       [4:0]    _zz_when_ArraySlice_l166_221_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_221_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_221_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_221_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_221;
  wire       [6:0]    _zz_when_ArraySlice_l113_221;
  wire       [6:0]    _zz_when_ArraySlice_l113_221_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_221_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_221_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_221_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_221;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_221_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_221_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_221_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_221;
  wire       [6:0]    _zz_when_ArraySlice_l118_221_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_221_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_221_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_221_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_221_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_221_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_221_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_221_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_221_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_222;
  wire       [5:0]    _zz_when_ArraySlice_l165_222_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_222;
  wire       [4:0]    _zz_when_ArraySlice_l166_222_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_222_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_222_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_222_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_222;
  wire       [6:0]    _zz_when_ArraySlice_l113_222;
  wire       [6:0]    _zz_when_ArraySlice_l113_222_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_222_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_222_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_222_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_222;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_222_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_222_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_222_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_222;
  wire       [6:0]    _zz_when_ArraySlice_l118_222_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_222_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_222_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_222_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_222_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_222_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_222_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_222_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_222_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_223;
  wire       [5:0]    _zz_when_ArraySlice_l165_223_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_223;
  wire       [3:0]    _zz_when_ArraySlice_l166_223_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_223_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_223_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_223_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_223;
  wire       [6:0]    _zz_when_ArraySlice_l113_223;
  wire       [6:0]    _zz_when_ArraySlice_l113_223_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_223_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_223_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_223_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_223;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_223_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_223_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_223_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_223;
  wire       [6:0]    _zz_when_ArraySlice_l118_223_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_223_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_223_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_223_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_223_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_223_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_223_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_223_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_223_8;
  wire                _zz_when_ArraySlice_l285;
  wire                _zz_when_ArraySlice_l285_1;
  wire                _zz_when_ArraySlice_l285_2;
  wire                _zz_when_ArraySlice_l285_3;
  wire                _zz_when_ArraySlice_l285_4;
  wire                _zz_when_ArraySlice_l285_5;
  wire       [5:0]    _zz_when_ArraySlice_l288;
  wire       [5:0]    _zz_when_ArraySlice_l288_1;
  wire       [5:0]    _zz_when_ArraySlice_l288_2;
  wire       [5:0]    _zz_when_ArraySlice_l288_3;
  wire       [5:0]    _zz_when_ArraySlice_l288_4;
  wire       [0:0]    _zz_when_ArraySlice_l288_5;
  wire       [5:0]    _zz_when_ArraySlice_l288_6;
  wire       [2:0]    _zz_when_ArraySlice_l288_7;
  wire       [5:0]    _zz_selectReadFifo_0_56;
  wire       [0:0]    _zz_selectReadFifo_0_57;
  wire       [12:0]   _zz_when_ArraySlice_l292;
  wire       [12:0]   _zz_when_ArraySlice_l292_1;
  wire       [12:0]   _zz_when_ArraySlice_l292_2;
  wire       [0:0]    _zz_when_ArraySlice_l292_3;
  wire       [12:0]   _zz_when_ArraySlice_l303;
  wire       [5:0]    _zz_when_ArraySlice_l303_1;
  wire       [5:0]    _zz_when_ArraySlice_l303_2;
  wire       [5:0]    _zz_when_ArraySlice_l303_3;
  wire       [0:0]    _zz_when_ArraySlice_l303_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_26;
  wire       [6:0]    _zz_when_ArraySlice_l95_26;
  wire       [6:0]    _zz_when_ArraySlice_l95_26_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_26_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_26_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_26_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_26;
  wire       [6:0]    _zz_when_ArraySlice_l99_26_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_8;
  wire       [6:0]    _zz_when_ArraySlice_l304_9;
  wire       [0:0]    _zz_when_ArraySlice_l304_10;
  wire       [6:0]    _zz_when_ArraySlice_l304_11;
  wire       [5:0]    _zz_selectReadFifo_0_58;
  wire       [5:0]    _zz_selectReadFifo_0_59;
  wire       [5:0]    _zz_selectReadFifo_0_60;
  wire       [0:0]    _zz_selectReadFifo_0_61;
  wire       [5:0]    _zz_when_ArraySlice_l165_224;
  wire       [5:0]    _zz_when_ArraySlice_l165_224_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_224_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_224;
  wire       [6:0]    _zz_when_ArraySlice_l166_224_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_224_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_224_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_224_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_224_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_224;
  wire       [6:0]    _zz_when_ArraySlice_l113_224;
  wire       [6:0]    _zz_when_ArraySlice_l113_224_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_224_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_224_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_224_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_224;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_224_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_224_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_224_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_224;
  wire       [6:0]    _zz_when_ArraySlice_l118_224_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_224_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_224_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_224_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_224_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_224_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_224_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_224_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_224_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_225;
  wire       [5:0]    _zz_when_ArraySlice_l165_225_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_225_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_225;
  wire       [5:0]    _zz_when_ArraySlice_l166_225_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_225_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_225_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_225_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_225;
  wire       [6:0]    _zz_when_ArraySlice_l113_225;
  wire       [6:0]    _zz_when_ArraySlice_l113_225_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_225_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_225_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_225_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_225;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_225_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_225_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_225_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_225;
  wire       [6:0]    _zz_when_ArraySlice_l118_225_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_225_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_225_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_225_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_225_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_225_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_225_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_225_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_225_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_225_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_226;
  wire       [5:0]    _zz_when_ArraySlice_l165_226_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_226_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_226;
  wire       [5:0]    _zz_when_ArraySlice_l166_226_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_226_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_226_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_226_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_226;
  wire       [6:0]    _zz_when_ArraySlice_l113_226;
  wire       [6:0]    _zz_when_ArraySlice_l113_226_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_226_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_226_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_226_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_226;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_226_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_226_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_226_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_226;
  wire       [6:0]    _zz_when_ArraySlice_l118_226_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_226_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_226_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_226_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_226_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_226_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_226_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_226_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_226_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_226_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_227;
  wire       [5:0]    _zz_when_ArraySlice_l165_227_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_227_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_227;
  wire       [5:0]    _zz_when_ArraySlice_l166_227_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_227_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_227_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_227_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_227;
  wire       [6:0]    _zz_when_ArraySlice_l113_227;
  wire       [6:0]    _zz_when_ArraySlice_l113_227_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_227_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_227_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_227_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_227;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_227_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_227_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_227_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_227;
  wire       [6:0]    _zz_when_ArraySlice_l118_227_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_227_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_227_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_227_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_227_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_227_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_227_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_227_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_227_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_227_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_228;
  wire       [5:0]    _zz_when_ArraySlice_l165_228_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_228;
  wire       [5:0]    _zz_when_ArraySlice_l166_228_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_228_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_228_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_228;
  wire       [6:0]    _zz_when_ArraySlice_l113_228;
  wire       [6:0]    _zz_when_ArraySlice_l113_228_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_228_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_228_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_228_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_228;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_228_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_228_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_228_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_228;
  wire       [6:0]    _zz_when_ArraySlice_l118_228_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_228_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_228_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_228_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_228_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_228_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_228_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_228_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_228_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_229;
  wire       [5:0]    _zz_when_ArraySlice_l165_229_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_229;
  wire       [4:0]    _zz_when_ArraySlice_l166_229_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_229_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_229_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_229_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_229;
  wire       [6:0]    _zz_when_ArraySlice_l113_229;
  wire       [6:0]    _zz_when_ArraySlice_l113_229_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_229_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_229_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_229_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_229;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_229_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_229_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_229_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_229;
  wire       [6:0]    _zz_when_ArraySlice_l118_229_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_229_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_229_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_229_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_229_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_229_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_229_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_229_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_229_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_230;
  wire       [5:0]    _zz_when_ArraySlice_l165_230_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_230;
  wire       [4:0]    _zz_when_ArraySlice_l166_230_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_230_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_230_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_230_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_230;
  wire       [6:0]    _zz_when_ArraySlice_l113_230;
  wire       [6:0]    _zz_when_ArraySlice_l113_230_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_230_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_230_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_230_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_230;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_230_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_230_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_230_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_230;
  wire       [6:0]    _zz_when_ArraySlice_l118_230_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_230_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_230_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_230_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_230_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_230_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_230_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_230_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_230_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_231;
  wire       [5:0]    _zz_when_ArraySlice_l165_231_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_231;
  wire       [3:0]    _zz_when_ArraySlice_l166_231_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_231_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_231_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_231_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_231;
  wire       [6:0]    _zz_when_ArraySlice_l113_231;
  wire       [6:0]    _zz_when_ArraySlice_l113_231_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_231_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_231_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_231_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_231;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_231_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_231_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_231_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_231;
  wire       [6:0]    _zz_when_ArraySlice_l118_231_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_231_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_231_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_231_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_231_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_231_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_231_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_231_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_231_8;
  wire                _zz_when_ArraySlice_l311;
  wire                _zz_when_ArraySlice_l311_1;
  wire                _zz_when_ArraySlice_l311_2;
  wire                _zz_when_ArraySlice_l311_3;
  wire                _zz_when_ArraySlice_l311_4;
  wire                _zz_when_ArraySlice_l311_5;
  wire       [5:0]    _zz_selectReadFifo_0_62;
  wire       [0:0]    _zz_selectReadFifo_0_63;
  wire       [12:0]   _zz_when_ArraySlice_l315;
  wire       [12:0]   _zz_when_ArraySlice_l315_1;
  wire       [12:0]   _zz_when_ArraySlice_l315_2;
  wire       [0:0]    _zz_when_ArraySlice_l315_3;
  wire       [5:0]    _zz_when_ArraySlice_l301;
  wire       [5:0]    _zz_when_ArraySlice_l301_1;
  wire       [2:0]    _zz_when_ArraySlice_l301_2;
  wire       [12:0]   _zz_when_ArraySlice_l322;
  wire       [5:0]    _zz_when_ArraySlice_l322_1;
  wire       [5:0]    _zz_when_ArraySlice_l322_2;
  wire       [5:0]    _zz_when_ArraySlice_l322_3;
  wire       [0:0]    _zz_when_ArraySlice_l322_4;
  wire       [5:0]    _zz_when_ArraySlice_l240_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l240_1_2;
  wire       [3:0]    _zz_when_ArraySlice_l240_1_3;
  reg        [6:0]    _zz_when_ArraySlice_l241_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l241_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l241_1_3;
  wire       [3:0]    _zz_when_ArraySlice_l241_1_4;
  wire       [5:0]    _zz__zz_outputStreamArrayData_1_valid_1_1;
  wire       [3:0]    _zz__zz_outputStreamArrayData_1_valid_1_2;
  reg                 _zz_outputStreamArrayData_1_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_1_payload_1;
  wire       [6:0]    _zz_when_ArraySlice_l247_1_1;
  wire       [0:0]    _zz_when_ArraySlice_l247_1_2;
  reg        [6:0]    _zz_when_ArraySlice_l247_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l247_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l247_1_5;
  wire       [3:0]    _zz_when_ArraySlice_l247_1_6;
  wire       [12:0]   _zz_when_ArraySlice_l248_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l248_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l248_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l248_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l248_1_5;
  wire       [5:0]    _zz_selectReadFifo_1_32;
  wire       [5:0]    _zz_selectReadFifo_1_33;
  wire       [5:0]    _zz_selectReadFifo_1_34;
  wire       [0:0]    _zz_selectReadFifo_1_35;
  wire       [5:0]    _zz_selectReadFifo_1_36;
  wire       [0:0]    _zz_selectReadFifo_1_37;
  wire       [12:0]   _zz_when_ArraySlice_l251_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l251_1_2;
  wire       [12:0]   _zz_when_ArraySlice_l251_1_3;
  wire       [0:0]    _zz_when_ArraySlice_l251_1_4;
  reg        [6:0]    _zz_when_ArraySlice_l256_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l256_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l256_1_3;
  wire       [3:0]    _zz_when_ArraySlice_l256_1_4;
  wire       [6:0]    _zz_when_ArraySlice_l256_1_5;
  wire       [0:0]    _zz_when_ArraySlice_l256_1_6;
  wire       [12:0]   _zz_when_ArraySlice_l257_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l257_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l257_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l257_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l257_1_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_27;
  wire       [6:0]    _zz_when_ArraySlice_l95_27;
  wire       [6:0]    _zz_when_ArraySlice_l95_27_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_27_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_27_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_27_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_1_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_1_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_1_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_27;
  wire       [6:0]    _zz_when_ArraySlice_l99_27_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_1_2;
  wire       [0:0]    _zz_when_ArraySlice_l259_1_3;
  wire       [6:0]    _zz_when_ArraySlice_l259_1_4;
  wire       [5:0]    _zz_selectReadFifo_1_38;
  wire       [5:0]    _zz_selectReadFifo_1_39;
  wire       [5:0]    _zz_selectReadFifo_1_40;
  wire       [0:0]    _zz_selectReadFifo_1_41;
  wire       [5:0]    _zz_selectReadFifo_1_42;
  wire       [5:0]    _zz_selectReadFifo_1_43;
  wire       [5:0]    _zz_selectReadFifo_1_44;
  wire       [0:0]    _zz_selectReadFifo_1_45;
  wire       [5:0]    _zz_when_ArraySlice_l165_232;
  wire       [5:0]    _zz_when_ArraySlice_l165_232_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_232_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_232;
  wire       [6:0]    _zz_when_ArraySlice_l166_232_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_232_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_232_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_232_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_232_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_232;
  wire       [6:0]    _zz_when_ArraySlice_l113_232;
  wire       [6:0]    _zz_when_ArraySlice_l113_232_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_232_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_232_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_232_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_232;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_232_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_232_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_232_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_232;
  wire       [6:0]    _zz_when_ArraySlice_l118_232_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_232_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_232_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_232_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_232_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_232_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_232_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_232_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_232_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_233;
  wire       [5:0]    _zz_when_ArraySlice_l165_233_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_233_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_233;
  wire       [5:0]    _zz_when_ArraySlice_l166_233_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_233_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_233_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_233_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_233;
  wire       [6:0]    _zz_when_ArraySlice_l113_233;
  wire       [6:0]    _zz_when_ArraySlice_l113_233_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_233_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_233_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_233_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_233;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_233_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_233_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_233_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_233;
  wire       [6:0]    _zz_when_ArraySlice_l118_233_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_233_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_233_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_233_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_233_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_233_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_233_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_233_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_233_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_233_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_234;
  wire       [5:0]    _zz_when_ArraySlice_l165_234_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_234_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_234;
  wire       [5:0]    _zz_when_ArraySlice_l166_234_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_234_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_234_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_234_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_234;
  wire       [6:0]    _zz_when_ArraySlice_l113_234;
  wire       [6:0]    _zz_when_ArraySlice_l113_234_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_234_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_234_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_234_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_234;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_234_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_234_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_234_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_234;
  wire       [6:0]    _zz_when_ArraySlice_l118_234_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_234_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_234_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_234_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_234_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_234_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_234_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_234_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_234_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_234_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_235;
  wire       [5:0]    _zz_when_ArraySlice_l165_235_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_235_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_235;
  wire       [5:0]    _zz_when_ArraySlice_l166_235_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_235_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_235_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_235_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_235;
  wire       [6:0]    _zz_when_ArraySlice_l113_235;
  wire       [6:0]    _zz_when_ArraySlice_l113_235_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_235_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_235_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_235_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_235;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_235_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_235_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_235_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_235;
  wire       [6:0]    _zz_when_ArraySlice_l118_235_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_235_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_235_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_235_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_235_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_235_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_235_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_235_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_235_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_235_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_236;
  wire       [5:0]    _zz_when_ArraySlice_l165_236_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_236;
  wire       [5:0]    _zz_when_ArraySlice_l166_236_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_236_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_236_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_236;
  wire       [6:0]    _zz_when_ArraySlice_l113_236;
  wire       [6:0]    _zz_when_ArraySlice_l113_236_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_236_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_236_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_236_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_236;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_236_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_236_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_236_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_236;
  wire       [6:0]    _zz_when_ArraySlice_l118_236_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_236_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_236_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_236_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_236_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_236_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_236_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_236_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_236_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_237;
  wire       [5:0]    _zz_when_ArraySlice_l165_237_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_237;
  wire       [4:0]    _zz_when_ArraySlice_l166_237_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_237_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_237_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_237_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_237;
  wire       [6:0]    _zz_when_ArraySlice_l113_237;
  wire       [6:0]    _zz_when_ArraySlice_l113_237_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_237_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_237_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_237_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_237;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_237_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_237_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_237_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_237;
  wire       [6:0]    _zz_when_ArraySlice_l118_237_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_237_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_237_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_237_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_237_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_237_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_237_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_237_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_237_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_238;
  wire       [5:0]    _zz_when_ArraySlice_l165_238_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_238;
  wire       [4:0]    _zz_when_ArraySlice_l166_238_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_238_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_238_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_238_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_238;
  wire       [6:0]    _zz_when_ArraySlice_l113_238;
  wire       [6:0]    _zz_when_ArraySlice_l113_238_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_238_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_238_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_238_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_238;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_238_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_238_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_238_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_238;
  wire       [6:0]    _zz_when_ArraySlice_l118_238_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_238_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_238_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_238_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_238_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_238_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_238_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_238_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_238_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_239;
  wire       [5:0]    _zz_when_ArraySlice_l165_239_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_239;
  wire       [3:0]    _zz_when_ArraySlice_l166_239_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_239_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_239_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_239_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_239;
  wire       [6:0]    _zz_when_ArraySlice_l113_239;
  wire       [6:0]    _zz_when_ArraySlice_l113_239_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_239_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_239_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_239_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_239;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_239_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_239_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_239_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_239;
  wire       [6:0]    _zz_when_ArraySlice_l118_239_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_239_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_239_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_239_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_239_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_239_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_239_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_239_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_239_8;
  wire                _zz_when_ArraySlice_l265_1_1;
  wire                _zz_when_ArraySlice_l265_1_2;
  wire                _zz_when_ArraySlice_l265_1_3;
  wire                _zz_when_ArraySlice_l265_1_4;
  wire                _zz_when_ArraySlice_l265_1_5;
  wire                _zz_when_ArraySlice_l265_1_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l268_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l268_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l268_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l268_1_5;
  wire       [0:0]    _zz_when_ArraySlice_l268_1_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_1_7;
  wire       [3:0]    _zz_when_ArraySlice_l268_1_8;
  wire       [5:0]    _zz_selectReadFifo_1_46;
  wire       [0:0]    _zz_selectReadFifo_1_47;
  wire       [12:0]   _zz_when_ArraySlice_l272_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l272_1_2;
  wire       [12:0]   _zz_when_ArraySlice_l272_1_3;
  wire       [0:0]    _zz_when_ArraySlice_l272_1_4;
  reg        [6:0]    _zz_when_ArraySlice_l276_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l276_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l276_1_3;
  wire       [3:0]    _zz_when_ArraySlice_l276_1_4;
  wire       [12:0]   _zz_when_ArraySlice_l277_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l277_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l277_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l277_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l277_1_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_28;
  wire       [6:0]    _zz_when_ArraySlice_l95_28;
  wire       [6:0]    _zz_when_ArraySlice_l95_28_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_28_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_28_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_28_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_1_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_1_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_1_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_28;
  wire       [6:0]    _zz_when_ArraySlice_l99_28_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_1_2;
  wire       [0:0]    _zz_when_ArraySlice_l279_1_3;
  wire       [6:0]    _zz_when_ArraySlice_l279_1_4;
  wire       [5:0]    _zz_selectReadFifo_1_48;
  wire       [5:0]    _zz_selectReadFifo_1_49;
  wire       [5:0]    _zz_selectReadFifo_1_50;
  wire       [0:0]    _zz_selectReadFifo_1_51;
  wire       [5:0]    _zz_selectReadFifo_1_52;
  wire       [5:0]    _zz_selectReadFifo_1_53;
  wire       [5:0]    _zz_selectReadFifo_1_54;
  wire       [0:0]    _zz_selectReadFifo_1_55;
  wire       [5:0]    _zz_when_ArraySlice_l165_240;
  wire       [5:0]    _zz_when_ArraySlice_l165_240_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_240_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_240;
  wire       [6:0]    _zz_when_ArraySlice_l166_240_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_240_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_240_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_240_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_240_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_240;
  wire       [6:0]    _zz_when_ArraySlice_l113_240;
  wire       [6:0]    _zz_when_ArraySlice_l113_240_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_240_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_240_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_240_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_240;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_240_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_240_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_240_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_240;
  wire       [6:0]    _zz_when_ArraySlice_l118_240_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_240_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_240_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_240_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_240_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_240_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_240_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_240_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_240_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_241;
  wire       [5:0]    _zz_when_ArraySlice_l165_241_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_241_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_241;
  wire       [5:0]    _zz_when_ArraySlice_l166_241_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_241_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_241_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_241_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_241;
  wire       [6:0]    _zz_when_ArraySlice_l113_241;
  wire       [6:0]    _zz_when_ArraySlice_l113_241_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_241_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_241_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_241_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_241;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_241_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_241_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_241_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_241;
  wire       [6:0]    _zz_when_ArraySlice_l118_241_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_241_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_241_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_241_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_241_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_241_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_241_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_241_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_241_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_241_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_242;
  wire       [5:0]    _zz_when_ArraySlice_l165_242_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_242_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_242;
  wire       [5:0]    _zz_when_ArraySlice_l166_242_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_242_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_242_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_242_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_242;
  wire       [6:0]    _zz_when_ArraySlice_l113_242;
  wire       [6:0]    _zz_when_ArraySlice_l113_242_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_242_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_242_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_242_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_242;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_242_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_242_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_242_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_242;
  wire       [6:0]    _zz_when_ArraySlice_l118_242_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_242_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_242_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_242_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_242_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_242_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_242_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_242_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_242_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_242_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_243;
  wire       [5:0]    _zz_when_ArraySlice_l165_243_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_243_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_243;
  wire       [5:0]    _zz_when_ArraySlice_l166_243_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_243_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_243_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_243_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_243;
  wire       [6:0]    _zz_when_ArraySlice_l113_243;
  wire       [6:0]    _zz_when_ArraySlice_l113_243_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_243_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_243_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_243_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_243;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_243_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_243_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_243_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_243;
  wire       [6:0]    _zz_when_ArraySlice_l118_243_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_243_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_243_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_243_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_243_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_243_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_243_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_243_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_243_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_243_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_244;
  wire       [5:0]    _zz_when_ArraySlice_l165_244_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_244;
  wire       [5:0]    _zz_when_ArraySlice_l166_244_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_244_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_244_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_244;
  wire       [6:0]    _zz_when_ArraySlice_l113_244;
  wire       [6:0]    _zz_when_ArraySlice_l113_244_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_244_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_244_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_244_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_244;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_244_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_244_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_244_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_244;
  wire       [6:0]    _zz_when_ArraySlice_l118_244_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_244_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_244_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_244_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_244_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_244_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_244_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_244_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_244_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_245;
  wire       [5:0]    _zz_when_ArraySlice_l165_245_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_245;
  wire       [4:0]    _zz_when_ArraySlice_l166_245_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_245_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_245_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_245_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_245;
  wire       [6:0]    _zz_when_ArraySlice_l113_245;
  wire       [6:0]    _zz_when_ArraySlice_l113_245_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_245_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_245_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_245_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_245;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_245_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_245_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_245_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_245;
  wire       [6:0]    _zz_when_ArraySlice_l118_245_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_245_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_245_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_245_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_245_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_245_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_245_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_245_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_245_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_246;
  wire       [5:0]    _zz_when_ArraySlice_l165_246_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_246;
  wire       [4:0]    _zz_when_ArraySlice_l166_246_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_246_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_246_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_246_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_246;
  wire       [6:0]    _zz_when_ArraySlice_l113_246;
  wire       [6:0]    _zz_when_ArraySlice_l113_246_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_246_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_246_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_246_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_246;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_246_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_246_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_246_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_246;
  wire       [6:0]    _zz_when_ArraySlice_l118_246_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_246_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_246_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_246_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_246_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_246_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_246_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_246_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_246_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_247;
  wire       [5:0]    _zz_when_ArraySlice_l165_247_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_247;
  wire       [3:0]    _zz_when_ArraySlice_l166_247_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_247_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_247_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_247_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_247;
  wire       [6:0]    _zz_when_ArraySlice_l113_247;
  wire       [6:0]    _zz_when_ArraySlice_l113_247_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_247_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_247_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_247_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_247;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_247_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_247_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_247_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_247;
  wire       [6:0]    _zz_when_ArraySlice_l118_247_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_247_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_247_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_247_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_247_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_247_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_247_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_247_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_247_8;
  wire                _zz_when_ArraySlice_l285_1_1;
  wire                _zz_when_ArraySlice_l285_1_2;
  wire                _zz_when_ArraySlice_l285_1_3;
  wire                _zz_when_ArraySlice_l285_1_4;
  wire                _zz_when_ArraySlice_l285_1_5;
  wire                _zz_when_ArraySlice_l285_1_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l288_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l288_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l288_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l288_1_5;
  wire       [0:0]    _zz_when_ArraySlice_l288_1_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_1_7;
  wire       [3:0]    _zz_when_ArraySlice_l288_1_8;
  wire       [5:0]    _zz_selectReadFifo_1_56;
  wire       [0:0]    _zz_selectReadFifo_1_57;
  wire       [12:0]   _zz_when_ArraySlice_l292_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l292_1_2;
  wire       [12:0]   _zz_when_ArraySlice_l292_1_3;
  wire       [0:0]    _zz_when_ArraySlice_l292_1_4;
  wire       [12:0]   _zz_when_ArraySlice_l303_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l303_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l303_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l303_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l303_1_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_29;
  wire       [6:0]    _zz_when_ArraySlice_l95_29;
  wire       [6:0]    _zz_when_ArraySlice_l95_29_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_29_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_29_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_29_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_1_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_1_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_1_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_29;
  wire       [6:0]    _zz_when_ArraySlice_l99_29_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_1_2;
  wire       [0:0]    _zz_when_ArraySlice_l304_1_3;
  wire       [6:0]    _zz_when_ArraySlice_l304_1_4;
  wire       [5:0]    _zz_selectReadFifo_1_58;
  wire       [5:0]    _zz_selectReadFifo_1_59;
  wire       [5:0]    _zz_selectReadFifo_1_60;
  wire       [0:0]    _zz_selectReadFifo_1_61;
  wire       [5:0]    _zz_when_ArraySlice_l165_248;
  wire       [5:0]    _zz_when_ArraySlice_l165_248_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_248_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_248;
  wire       [6:0]    _zz_when_ArraySlice_l166_248_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_248_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_248_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_248_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_248_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_248;
  wire       [6:0]    _zz_when_ArraySlice_l113_248;
  wire       [6:0]    _zz_when_ArraySlice_l113_248_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_248_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_248_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_248_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_248;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_248_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_248_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_248_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_248;
  wire       [6:0]    _zz_when_ArraySlice_l118_248_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_248_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_248_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_248_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_248_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_248_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_248_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_248_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_248_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_249;
  wire       [5:0]    _zz_when_ArraySlice_l165_249_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_249_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_249;
  wire       [5:0]    _zz_when_ArraySlice_l166_249_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_249_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_249_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_249_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_249;
  wire       [6:0]    _zz_when_ArraySlice_l113_249;
  wire       [6:0]    _zz_when_ArraySlice_l113_249_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_249_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_249_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_249_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_249;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_249_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_249_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_249_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_249;
  wire       [6:0]    _zz_when_ArraySlice_l118_249_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_249_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_249_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_249_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_249_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_249_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_249_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_249_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_249_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_249_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_250;
  wire       [5:0]    _zz_when_ArraySlice_l165_250_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_250_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_250;
  wire       [5:0]    _zz_when_ArraySlice_l166_250_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_250_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_250_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_250_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_250;
  wire       [6:0]    _zz_when_ArraySlice_l113_250;
  wire       [6:0]    _zz_when_ArraySlice_l113_250_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_250_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_250_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_250_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_250;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_250_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_250_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_250_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_250;
  wire       [6:0]    _zz_when_ArraySlice_l118_250_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_250_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_250_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_250_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_250_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_250_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_250_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_250_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_250_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_250_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_251;
  wire       [5:0]    _zz_when_ArraySlice_l165_251_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_251_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_251;
  wire       [5:0]    _zz_when_ArraySlice_l166_251_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_251_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_251_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_251_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_251;
  wire       [6:0]    _zz_when_ArraySlice_l113_251;
  wire       [6:0]    _zz_when_ArraySlice_l113_251_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_251_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_251_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_251_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_251;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_251_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_251_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_251_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_251;
  wire       [6:0]    _zz_when_ArraySlice_l118_251_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_251_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_251_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_251_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_251_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_251_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_251_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_251_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_251_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_251_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_252;
  wire       [5:0]    _zz_when_ArraySlice_l165_252_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_252;
  wire       [5:0]    _zz_when_ArraySlice_l166_252_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_252_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_252_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_252;
  wire       [6:0]    _zz_when_ArraySlice_l113_252;
  wire       [6:0]    _zz_when_ArraySlice_l113_252_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_252_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_252_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_252_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_252;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_252_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_252_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_252_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_252;
  wire       [6:0]    _zz_when_ArraySlice_l118_252_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_252_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_252_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_252_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_252_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_252_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_252_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_252_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_252_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_253;
  wire       [5:0]    _zz_when_ArraySlice_l165_253_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_253;
  wire       [4:0]    _zz_when_ArraySlice_l166_253_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_253_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_253_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_253_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_253;
  wire       [6:0]    _zz_when_ArraySlice_l113_253;
  wire       [6:0]    _zz_when_ArraySlice_l113_253_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_253_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_253_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_253_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_253;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_253_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_253_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_253_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_253;
  wire       [6:0]    _zz_when_ArraySlice_l118_253_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_253_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_253_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_253_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_253_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_253_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_253_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_253_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_253_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_254;
  wire       [5:0]    _zz_when_ArraySlice_l165_254_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_254;
  wire       [4:0]    _zz_when_ArraySlice_l166_254_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_254_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_254_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_254_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_254;
  wire       [6:0]    _zz_when_ArraySlice_l113_254;
  wire       [6:0]    _zz_when_ArraySlice_l113_254_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_254_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_254_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_254_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_254;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_254_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_254_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_254_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_254;
  wire       [6:0]    _zz_when_ArraySlice_l118_254_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_254_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_254_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_254_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_254_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_254_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_254_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_254_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_254_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_255;
  wire       [5:0]    _zz_when_ArraySlice_l165_255_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_255;
  wire       [3:0]    _zz_when_ArraySlice_l166_255_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_255_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_255_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_255_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_255;
  wire       [6:0]    _zz_when_ArraySlice_l113_255;
  wire       [6:0]    _zz_when_ArraySlice_l113_255_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_255_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_255_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_255_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_255;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_255_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_255_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_255_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_255;
  wire       [6:0]    _zz_when_ArraySlice_l118_255_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_255_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_255_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_255_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_255_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_255_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_255_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_255_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_255_8;
  wire                _zz_when_ArraySlice_l311_1_1;
  wire                _zz_when_ArraySlice_l311_1_2;
  wire                _zz_when_ArraySlice_l311_1_3;
  wire                _zz_when_ArraySlice_l311_1_4;
  wire                _zz_when_ArraySlice_l311_1_5;
  wire                _zz_when_ArraySlice_l311_1_6;
  wire       [5:0]    _zz_selectReadFifo_1_62;
  wire       [0:0]    _zz_selectReadFifo_1_63;
  wire       [12:0]   _zz_when_ArraySlice_l315_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l315_1_2;
  wire       [12:0]   _zz_when_ArraySlice_l315_1_3;
  wire       [0:0]    _zz_when_ArraySlice_l315_1_4;
  wire       [5:0]    _zz_when_ArraySlice_l301_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l301_1_2;
  wire       [3:0]    _zz_when_ArraySlice_l301_1_3;
  wire       [12:0]   _zz_when_ArraySlice_l322_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l322_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l322_1_3;
  wire       [5:0]    _zz_when_ArraySlice_l322_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l322_1_5;
  wire       [5:0]    _zz_when_ArraySlice_l240_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l240_2_2;
  wire       [4:0]    _zz_when_ArraySlice_l240_2_3;
  reg        [6:0]    _zz_when_ArraySlice_l241_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l241_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l241_2_3;
  wire       [4:0]    _zz_when_ArraySlice_l241_2_4;
  wire       [5:0]    _zz__zz_outputStreamArrayData_2_valid_1_1;
  wire       [4:0]    _zz__zz_outputStreamArrayData_2_valid_1_2;
  reg                 _zz_outputStreamArrayData_2_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_2_payload_1;
  wire       [6:0]    _zz_when_ArraySlice_l247_2_1;
  wire       [0:0]    _zz_when_ArraySlice_l247_2_2;
  reg        [6:0]    _zz_when_ArraySlice_l247_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l247_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l247_2_5;
  wire       [4:0]    _zz_when_ArraySlice_l247_2_6;
  wire       [12:0]   _zz_when_ArraySlice_l248_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l248_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l248_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l248_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l248_2_5;
  wire       [5:0]    _zz_selectReadFifo_2_32;
  wire       [5:0]    _zz_selectReadFifo_2_33;
  wire       [5:0]    _zz_selectReadFifo_2_34;
  wire       [0:0]    _zz_selectReadFifo_2_35;
  wire       [5:0]    _zz_selectReadFifo_2_36;
  wire       [0:0]    _zz_selectReadFifo_2_37;
  wire       [12:0]   _zz_when_ArraySlice_l251_2_1;
  wire       [12:0]   _zz_when_ArraySlice_l251_2_2;
  wire       [12:0]   _zz_when_ArraySlice_l251_2_3;
  wire       [0:0]    _zz_when_ArraySlice_l251_2_4;
  reg        [6:0]    _zz_when_ArraySlice_l256_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l256_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l256_2_3;
  wire       [4:0]    _zz_when_ArraySlice_l256_2_4;
  wire       [6:0]    _zz_when_ArraySlice_l256_2_5;
  wire       [0:0]    _zz_when_ArraySlice_l256_2_6;
  wire       [12:0]   _zz_when_ArraySlice_l257_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l257_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l257_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l257_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l257_2_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_30;
  wire       [6:0]    _zz_when_ArraySlice_l95_30;
  wire       [6:0]    _zz_when_ArraySlice_l95_30_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_30_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_30_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_30_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_2_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_2_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_2_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_30;
  wire       [6:0]    _zz_when_ArraySlice_l99_30_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_2_2;
  wire       [0:0]    _zz_when_ArraySlice_l259_2_3;
  wire       [6:0]    _zz_when_ArraySlice_l259_2_4;
  wire       [5:0]    _zz_selectReadFifo_2_38;
  wire       [5:0]    _zz_selectReadFifo_2_39;
  wire       [5:0]    _zz_selectReadFifo_2_40;
  wire       [0:0]    _zz_selectReadFifo_2_41;
  wire       [5:0]    _zz_selectReadFifo_2_42;
  wire       [5:0]    _zz_selectReadFifo_2_43;
  wire       [5:0]    _zz_selectReadFifo_2_44;
  wire       [0:0]    _zz_selectReadFifo_2_45;
  wire       [5:0]    _zz_when_ArraySlice_l165_256;
  wire       [5:0]    _zz_when_ArraySlice_l165_256_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_256_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_256;
  wire       [6:0]    _zz_when_ArraySlice_l166_256_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_256_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_256_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_256_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_256_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_256;
  wire       [6:0]    _zz_when_ArraySlice_l113_256;
  wire       [6:0]    _zz_when_ArraySlice_l113_256_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_256_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_256_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_256_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_256;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_256_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_256_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_256_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_256;
  wire       [6:0]    _zz_when_ArraySlice_l118_256_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_256_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_256_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_256_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_256_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_256_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_256_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_256_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_256_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_257;
  wire       [5:0]    _zz_when_ArraySlice_l165_257_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_257_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_257;
  wire       [5:0]    _zz_when_ArraySlice_l166_257_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_257_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_257_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_257_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_257;
  wire       [6:0]    _zz_when_ArraySlice_l113_257;
  wire       [6:0]    _zz_when_ArraySlice_l113_257_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_257_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_257_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_257_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_257;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_257_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_257_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_257_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_257;
  wire       [6:0]    _zz_when_ArraySlice_l118_257_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_257_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_257_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_257_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_257_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_257_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_257_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_257_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_257_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_257_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_258;
  wire       [5:0]    _zz_when_ArraySlice_l165_258_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_258_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_258;
  wire       [5:0]    _zz_when_ArraySlice_l166_258_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_258_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_258_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_258_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_258;
  wire       [6:0]    _zz_when_ArraySlice_l113_258;
  wire       [6:0]    _zz_when_ArraySlice_l113_258_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_258_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_258_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_258_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_258;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_258_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_258_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_258_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_258;
  wire       [6:0]    _zz_when_ArraySlice_l118_258_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_258_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_258_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_258_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_258_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_258_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_258_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_258_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_258_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_258_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_259;
  wire       [5:0]    _zz_when_ArraySlice_l165_259_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_259_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_259;
  wire       [5:0]    _zz_when_ArraySlice_l166_259_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_259_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_259_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_259_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_259;
  wire       [6:0]    _zz_when_ArraySlice_l113_259;
  wire       [6:0]    _zz_when_ArraySlice_l113_259_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_259_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_259_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_259_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_259;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_259_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_259_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_259_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_259;
  wire       [6:0]    _zz_when_ArraySlice_l118_259_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_259_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_259_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_259_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_259_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_259_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_259_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_259_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_259_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_259_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_260;
  wire       [5:0]    _zz_when_ArraySlice_l165_260_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_260;
  wire       [5:0]    _zz_when_ArraySlice_l166_260_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_260_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_260_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_260;
  wire       [6:0]    _zz_when_ArraySlice_l113_260;
  wire       [6:0]    _zz_when_ArraySlice_l113_260_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_260_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_260_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_260_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_260;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_260_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_260_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_260_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_260;
  wire       [6:0]    _zz_when_ArraySlice_l118_260_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_260_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_260_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_260_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_260_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_260_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_260_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_260_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_260_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_261;
  wire       [5:0]    _zz_when_ArraySlice_l165_261_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_261;
  wire       [4:0]    _zz_when_ArraySlice_l166_261_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_261_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_261_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_261_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_261;
  wire       [6:0]    _zz_when_ArraySlice_l113_261;
  wire       [6:0]    _zz_when_ArraySlice_l113_261_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_261_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_261_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_261_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_261;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_261_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_261_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_261_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_261;
  wire       [6:0]    _zz_when_ArraySlice_l118_261_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_261_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_261_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_261_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_261_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_261_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_261_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_261_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_261_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_262;
  wire       [5:0]    _zz_when_ArraySlice_l165_262_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_262;
  wire       [4:0]    _zz_when_ArraySlice_l166_262_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_262_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_262_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_262_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_262;
  wire       [6:0]    _zz_when_ArraySlice_l113_262;
  wire       [6:0]    _zz_when_ArraySlice_l113_262_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_262_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_262_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_262_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_262;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_262_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_262_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_262_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_262;
  wire       [6:0]    _zz_when_ArraySlice_l118_262_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_262_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_262_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_262_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_262_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_262_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_262_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_262_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_262_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_263;
  wire       [5:0]    _zz_when_ArraySlice_l165_263_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_263;
  wire       [3:0]    _zz_when_ArraySlice_l166_263_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_263_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_263_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_263_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_263;
  wire       [6:0]    _zz_when_ArraySlice_l113_263;
  wire       [6:0]    _zz_when_ArraySlice_l113_263_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_263_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_263_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_263_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_263;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_263_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_263_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_263_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_263;
  wire       [6:0]    _zz_when_ArraySlice_l118_263_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_263_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_263_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_263_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_263_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_263_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_263_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_263_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_263_8;
  wire                _zz_when_ArraySlice_l265_2_1;
  wire                _zz_when_ArraySlice_l265_2_2;
  wire                _zz_when_ArraySlice_l265_2_3;
  wire                _zz_when_ArraySlice_l265_2_4;
  wire                _zz_when_ArraySlice_l265_2_5;
  wire                _zz_when_ArraySlice_l265_2_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l268_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l268_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l268_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l268_2_5;
  wire       [0:0]    _zz_when_ArraySlice_l268_2_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_2_7;
  wire       [4:0]    _zz_when_ArraySlice_l268_2_8;
  wire       [5:0]    _zz_selectReadFifo_2_46;
  wire       [0:0]    _zz_selectReadFifo_2_47;
  wire       [12:0]   _zz_when_ArraySlice_l272_2_1;
  wire       [12:0]   _zz_when_ArraySlice_l272_2_2;
  wire       [12:0]   _zz_when_ArraySlice_l272_2_3;
  wire       [0:0]    _zz_when_ArraySlice_l272_2_4;
  reg        [6:0]    _zz_when_ArraySlice_l276_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l276_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l276_2_3;
  wire       [4:0]    _zz_when_ArraySlice_l276_2_4;
  wire       [12:0]   _zz_when_ArraySlice_l277_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l277_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l277_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l277_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l277_2_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_31;
  wire       [6:0]    _zz_when_ArraySlice_l95_31;
  wire       [6:0]    _zz_when_ArraySlice_l95_31_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_31_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_31_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_31_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_2_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_2_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_2_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_31;
  wire       [6:0]    _zz_when_ArraySlice_l99_31_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_2_2;
  wire       [0:0]    _zz_when_ArraySlice_l279_2_3;
  wire       [6:0]    _zz_when_ArraySlice_l279_2_4;
  wire       [5:0]    _zz_selectReadFifo_2_48;
  wire       [5:0]    _zz_selectReadFifo_2_49;
  wire       [5:0]    _zz_selectReadFifo_2_50;
  wire       [0:0]    _zz_selectReadFifo_2_51;
  wire       [5:0]    _zz_selectReadFifo_2_52;
  wire       [5:0]    _zz_selectReadFifo_2_53;
  wire       [5:0]    _zz_selectReadFifo_2_54;
  wire       [0:0]    _zz_selectReadFifo_2_55;
  wire       [5:0]    _zz_when_ArraySlice_l165_264;
  wire       [5:0]    _zz_when_ArraySlice_l165_264_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_264_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_264;
  wire       [6:0]    _zz_when_ArraySlice_l166_264_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_264_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_264_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_264_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_264_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_264;
  wire       [6:0]    _zz_when_ArraySlice_l113_264;
  wire       [6:0]    _zz_when_ArraySlice_l113_264_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_264_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_264_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_264_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_264;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_264_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_264_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_264_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_264;
  wire       [6:0]    _zz_when_ArraySlice_l118_264_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_264_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_264_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_264_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_264_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_264_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_264_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_264_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_264_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_265;
  wire       [5:0]    _zz_when_ArraySlice_l165_265_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_265_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_265;
  wire       [5:0]    _zz_when_ArraySlice_l166_265_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_265_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_265_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_265_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_265;
  wire       [6:0]    _zz_when_ArraySlice_l113_265;
  wire       [6:0]    _zz_when_ArraySlice_l113_265_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_265_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_265_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_265_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_265;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_265_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_265_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_265_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_265;
  wire       [6:0]    _zz_when_ArraySlice_l118_265_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_265_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_265_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_265_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_265_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_265_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_265_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_265_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_265_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_265_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_266;
  wire       [5:0]    _zz_when_ArraySlice_l165_266_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_266_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_266;
  wire       [5:0]    _zz_when_ArraySlice_l166_266_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_266_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_266_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_266_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_266;
  wire       [6:0]    _zz_when_ArraySlice_l113_266;
  wire       [6:0]    _zz_when_ArraySlice_l113_266_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_266_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_266_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_266_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_266;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_266_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_266_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_266_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_266;
  wire       [6:0]    _zz_when_ArraySlice_l118_266_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_266_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_266_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_266_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_266_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_266_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_266_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_266_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_266_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_266_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_267;
  wire       [5:0]    _zz_when_ArraySlice_l165_267_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_267_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_267;
  wire       [5:0]    _zz_when_ArraySlice_l166_267_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_267_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_267_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_267_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_267;
  wire       [6:0]    _zz_when_ArraySlice_l113_267;
  wire       [6:0]    _zz_when_ArraySlice_l113_267_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_267_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_267_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_267_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_267;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_267_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_267_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_267_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_267;
  wire       [6:0]    _zz_when_ArraySlice_l118_267_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_267_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_267_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_267_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_267_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_267_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_267_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_267_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_267_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_267_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_268;
  wire       [5:0]    _zz_when_ArraySlice_l165_268_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_268;
  wire       [5:0]    _zz_when_ArraySlice_l166_268_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_268_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_268_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_268;
  wire       [6:0]    _zz_when_ArraySlice_l113_268;
  wire       [6:0]    _zz_when_ArraySlice_l113_268_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_268_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_268_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_268_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_268;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_268_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_268_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_268_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_268;
  wire       [6:0]    _zz_when_ArraySlice_l118_268_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_268_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_268_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_268_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_268_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_268_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_268_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_268_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_268_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_269;
  wire       [5:0]    _zz_when_ArraySlice_l165_269_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_269;
  wire       [4:0]    _zz_when_ArraySlice_l166_269_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_269_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_269_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_269_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_269;
  wire       [6:0]    _zz_when_ArraySlice_l113_269;
  wire       [6:0]    _zz_when_ArraySlice_l113_269_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_269_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_269_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_269_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_269;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_269_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_269_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_269_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_269;
  wire       [6:0]    _zz_when_ArraySlice_l118_269_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_269_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_269_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_269_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_269_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_269_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_269_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_269_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_269_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_270;
  wire       [5:0]    _zz_when_ArraySlice_l165_270_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_270;
  wire       [4:0]    _zz_when_ArraySlice_l166_270_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_270_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_270_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_270_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_270;
  wire       [6:0]    _zz_when_ArraySlice_l113_270;
  wire       [6:0]    _zz_when_ArraySlice_l113_270_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_270_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_270_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_270_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_270;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_270_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_270_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_270_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_270;
  wire       [6:0]    _zz_when_ArraySlice_l118_270_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_270_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_270_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_270_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_270_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_270_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_270_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_270_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_270_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_271;
  wire       [5:0]    _zz_when_ArraySlice_l165_271_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_271;
  wire       [3:0]    _zz_when_ArraySlice_l166_271_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_271_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_271_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_271_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_271;
  wire       [6:0]    _zz_when_ArraySlice_l113_271;
  wire       [6:0]    _zz_when_ArraySlice_l113_271_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_271_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_271_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_271_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_271;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_271_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_271_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_271_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_271;
  wire       [6:0]    _zz_when_ArraySlice_l118_271_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_271_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_271_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_271_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_271_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_271_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_271_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_271_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_271_8;
  wire                _zz_when_ArraySlice_l285_2_1;
  wire                _zz_when_ArraySlice_l285_2_2;
  wire                _zz_when_ArraySlice_l285_2_3;
  wire                _zz_when_ArraySlice_l285_2_4;
  wire                _zz_when_ArraySlice_l285_2_5;
  wire                _zz_when_ArraySlice_l285_2_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l288_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l288_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l288_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l288_2_5;
  wire       [0:0]    _zz_when_ArraySlice_l288_2_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_2_7;
  wire       [4:0]    _zz_when_ArraySlice_l288_2_8;
  wire       [5:0]    _zz_selectReadFifo_2_56;
  wire       [0:0]    _zz_selectReadFifo_2_57;
  wire       [12:0]   _zz_when_ArraySlice_l292_2_1;
  wire       [12:0]   _zz_when_ArraySlice_l292_2_2;
  wire       [12:0]   _zz_when_ArraySlice_l292_2_3;
  wire       [0:0]    _zz_when_ArraySlice_l292_2_4;
  wire       [12:0]   _zz_when_ArraySlice_l303_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l303_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l303_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l303_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l303_2_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_32;
  wire       [6:0]    _zz_when_ArraySlice_l95_32;
  wire       [6:0]    _zz_when_ArraySlice_l95_32_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_32_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_32_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_32_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_2_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_2_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_2_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_32;
  wire       [6:0]    _zz_when_ArraySlice_l99_32_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_2_2;
  wire       [0:0]    _zz_when_ArraySlice_l304_2_3;
  wire       [6:0]    _zz_when_ArraySlice_l304_2_4;
  wire       [5:0]    _zz_selectReadFifo_2_58;
  wire       [5:0]    _zz_selectReadFifo_2_59;
  wire       [5:0]    _zz_selectReadFifo_2_60;
  wire       [0:0]    _zz_selectReadFifo_2_61;
  wire       [5:0]    _zz_when_ArraySlice_l165_272;
  wire       [5:0]    _zz_when_ArraySlice_l165_272_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_272_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_272;
  wire       [6:0]    _zz_when_ArraySlice_l166_272_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_272_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_272_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_272_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_272_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_272;
  wire       [6:0]    _zz_when_ArraySlice_l113_272;
  wire       [6:0]    _zz_when_ArraySlice_l113_272_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_272_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_272_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_272_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_272;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_272_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_272_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_272_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_272;
  wire       [6:0]    _zz_when_ArraySlice_l118_272_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_272_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_272_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_272_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_272_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_272_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_272_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_272_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_272_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_273;
  wire       [5:0]    _zz_when_ArraySlice_l165_273_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_273_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_273;
  wire       [5:0]    _zz_when_ArraySlice_l166_273_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_273_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_273_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_273_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_273;
  wire       [6:0]    _zz_when_ArraySlice_l113_273;
  wire       [6:0]    _zz_when_ArraySlice_l113_273_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_273_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_273_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_273_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_273;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_273_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_273_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_273_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_273;
  wire       [6:0]    _zz_when_ArraySlice_l118_273_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_273_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_273_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_273_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_273_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_273_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_273_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_273_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_273_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_273_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_274;
  wire       [5:0]    _zz_when_ArraySlice_l165_274_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_274_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_274;
  wire       [5:0]    _zz_when_ArraySlice_l166_274_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_274_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_274_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_274_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_274;
  wire       [6:0]    _zz_when_ArraySlice_l113_274;
  wire       [6:0]    _zz_when_ArraySlice_l113_274_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_274_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_274_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_274_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_274;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_274_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_274_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_274_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_274;
  wire       [6:0]    _zz_when_ArraySlice_l118_274_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_274_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_274_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_274_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_274_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_274_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_274_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_274_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_274_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_274_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_275;
  wire       [5:0]    _zz_when_ArraySlice_l165_275_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_275_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_275;
  wire       [5:0]    _zz_when_ArraySlice_l166_275_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_275_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_275_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_275_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_275;
  wire       [6:0]    _zz_when_ArraySlice_l113_275;
  wire       [6:0]    _zz_when_ArraySlice_l113_275_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_275_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_275_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_275_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_275;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_275_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_275_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_275_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_275;
  wire       [6:0]    _zz_when_ArraySlice_l118_275_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_275_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_275_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_275_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_275_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_275_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_275_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_275_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_275_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_275_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_276;
  wire       [5:0]    _zz_when_ArraySlice_l165_276_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_276;
  wire       [5:0]    _zz_when_ArraySlice_l166_276_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_276_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_276_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_276;
  wire       [6:0]    _zz_when_ArraySlice_l113_276;
  wire       [6:0]    _zz_when_ArraySlice_l113_276_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_276_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_276_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_276_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_276;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_276_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_276_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_276_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_276;
  wire       [6:0]    _zz_when_ArraySlice_l118_276_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_276_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_276_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_276_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_276_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_276_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_276_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_276_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_276_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_277;
  wire       [5:0]    _zz_when_ArraySlice_l165_277_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_277;
  wire       [4:0]    _zz_when_ArraySlice_l166_277_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_277_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_277_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_277_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_277;
  wire       [6:0]    _zz_when_ArraySlice_l113_277;
  wire       [6:0]    _zz_when_ArraySlice_l113_277_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_277_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_277_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_277_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_277;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_277_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_277_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_277_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_277;
  wire       [6:0]    _zz_when_ArraySlice_l118_277_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_277_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_277_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_277_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_277_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_277_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_277_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_277_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_277_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_278;
  wire       [5:0]    _zz_when_ArraySlice_l165_278_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_278;
  wire       [4:0]    _zz_when_ArraySlice_l166_278_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_278_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_278_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_278_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_278;
  wire       [6:0]    _zz_when_ArraySlice_l113_278;
  wire       [6:0]    _zz_when_ArraySlice_l113_278_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_278_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_278_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_278_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_278;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_278_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_278_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_278_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_278;
  wire       [6:0]    _zz_when_ArraySlice_l118_278_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_278_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_278_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_278_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_278_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_278_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_278_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_278_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_278_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_279;
  wire       [5:0]    _zz_when_ArraySlice_l165_279_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_279;
  wire       [3:0]    _zz_when_ArraySlice_l166_279_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_279_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_279_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_279_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_279;
  wire       [6:0]    _zz_when_ArraySlice_l113_279;
  wire       [6:0]    _zz_when_ArraySlice_l113_279_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_279_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_279_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_279_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_279;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_279_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_279_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_279_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_279;
  wire       [6:0]    _zz_when_ArraySlice_l118_279_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_279_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_279_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_279_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_279_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_279_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_279_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_279_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_279_8;
  wire                _zz_when_ArraySlice_l311_2_1;
  wire                _zz_when_ArraySlice_l311_2_2;
  wire                _zz_when_ArraySlice_l311_2_3;
  wire                _zz_when_ArraySlice_l311_2_4;
  wire                _zz_when_ArraySlice_l311_2_5;
  wire                _zz_when_ArraySlice_l311_2_6;
  wire       [5:0]    _zz_selectReadFifo_2_62;
  wire       [0:0]    _zz_selectReadFifo_2_63;
  wire       [12:0]   _zz_when_ArraySlice_l315_2_1;
  wire       [12:0]   _zz_when_ArraySlice_l315_2_2;
  wire       [12:0]   _zz_when_ArraySlice_l315_2_3;
  wire       [0:0]    _zz_when_ArraySlice_l315_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l301_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l301_2_2;
  wire       [4:0]    _zz_when_ArraySlice_l301_2_3;
  wire       [12:0]   _zz_when_ArraySlice_l322_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l322_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l322_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l322_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l322_2_5;
  wire       [5:0]    _zz_when_ArraySlice_l240_3;
  wire       [5:0]    _zz_when_ArraySlice_l240_3_1;
  wire       [4:0]    _zz_when_ArraySlice_l240_3_2;
  reg        [6:0]    _zz_when_ArraySlice_l241_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l241_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l241_3_3;
  wire       [4:0]    _zz_when_ArraySlice_l241_3_4;
  wire       [5:0]    _zz__zz_outputStreamArrayData_3_valid_1_1;
  wire       [4:0]    _zz__zz_outputStreamArrayData_3_valid_1_2;
  reg                 _zz_outputStreamArrayData_3_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_3_payload_1;
  wire       [6:0]    _zz_when_ArraySlice_l247_3_1;
  wire       [0:0]    _zz_when_ArraySlice_l247_3_2;
  reg        [6:0]    _zz_when_ArraySlice_l247_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l247_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l247_3_5;
  wire       [4:0]    _zz_when_ArraySlice_l247_3_6;
  wire       [12:0]   _zz_when_ArraySlice_l248_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l248_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l248_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l248_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l248_3_5;
  wire       [5:0]    _zz_selectReadFifo_3_32;
  wire       [5:0]    _zz_selectReadFifo_3_33;
  wire       [5:0]    _zz_selectReadFifo_3_34;
  wire       [0:0]    _zz_selectReadFifo_3_35;
  wire       [5:0]    _zz_selectReadFifo_3_36;
  wire       [0:0]    _zz_selectReadFifo_3_37;
  wire       [12:0]   _zz_when_ArraySlice_l251_3_1;
  wire       [12:0]   _zz_when_ArraySlice_l251_3_2;
  wire       [12:0]   _zz_when_ArraySlice_l251_3_3;
  wire       [0:0]    _zz_when_ArraySlice_l251_3_4;
  reg        [6:0]    _zz_when_ArraySlice_l256_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l256_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l256_3_3;
  wire       [4:0]    _zz_when_ArraySlice_l256_3_4;
  wire       [6:0]    _zz_when_ArraySlice_l256_3_5;
  wire       [0:0]    _zz_when_ArraySlice_l256_3_6;
  wire       [12:0]   _zz_when_ArraySlice_l257_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l257_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l257_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l257_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l257_3_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_33;
  wire       [6:0]    _zz_when_ArraySlice_l95_33;
  wire       [6:0]    _zz_when_ArraySlice_l95_33_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_33_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_33_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_33_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_3_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_3_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_3_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_33;
  wire       [6:0]    _zz_when_ArraySlice_l99_33_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_3_2;
  wire       [0:0]    _zz_when_ArraySlice_l259_3_3;
  wire       [6:0]    _zz_when_ArraySlice_l259_3_4;
  wire       [5:0]    _zz_selectReadFifo_3_38;
  wire       [5:0]    _zz_selectReadFifo_3_39;
  wire       [5:0]    _zz_selectReadFifo_3_40;
  wire       [0:0]    _zz_selectReadFifo_3_41;
  wire       [5:0]    _zz_selectReadFifo_3_42;
  wire       [5:0]    _zz_selectReadFifo_3_43;
  wire       [5:0]    _zz_selectReadFifo_3_44;
  wire       [0:0]    _zz_selectReadFifo_3_45;
  wire       [5:0]    _zz_when_ArraySlice_l165_280;
  wire       [5:0]    _zz_when_ArraySlice_l165_280_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_280_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_280;
  wire       [6:0]    _zz_when_ArraySlice_l166_280_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_280_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_280_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_280_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_280_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_280;
  wire       [6:0]    _zz_when_ArraySlice_l113_280;
  wire       [6:0]    _zz_when_ArraySlice_l113_280_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_280_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_280_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_280_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_280;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_280_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_280_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_280_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_280;
  wire       [6:0]    _zz_when_ArraySlice_l118_280_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_280_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_280_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_280_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_280_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_280_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_280_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_280_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_280_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_281;
  wire       [5:0]    _zz_when_ArraySlice_l165_281_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_281_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_281;
  wire       [5:0]    _zz_when_ArraySlice_l166_281_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_281_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_281_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_281_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_281;
  wire       [6:0]    _zz_when_ArraySlice_l113_281;
  wire       [6:0]    _zz_when_ArraySlice_l113_281_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_281_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_281_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_281_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_281;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_281_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_281_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_281_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_281;
  wire       [6:0]    _zz_when_ArraySlice_l118_281_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_281_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_281_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_281_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_281_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_281_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_281_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_281_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_281_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_281_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_282;
  wire       [5:0]    _zz_when_ArraySlice_l165_282_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_282_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_282;
  wire       [5:0]    _zz_when_ArraySlice_l166_282_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_282_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_282_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_282_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_282;
  wire       [6:0]    _zz_when_ArraySlice_l113_282;
  wire       [6:0]    _zz_when_ArraySlice_l113_282_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_282_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_282_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_282_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_282;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_282_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_282_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_282_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_282;
  wire       [6:0]    _zz_when_ArraySlice_l118_282_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_282_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_282_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_282_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_282_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_282_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_282_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_282_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_282_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_282_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_283;
  wire       [5:0]    _zz_when_ArraySlice_l165_283_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_283_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_283;
  wire       [5:0]    _zz_when_ArraySlice_l166_283_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_283_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_283_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_283_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_283;
  wire       [6:0]    _zz_when_ArraySlice_l113_283;
  wire       [6:0]    _zz_when_ArraySlice_l113_283_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_283_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_283_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_283_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_283;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_283_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_283_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_283_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_283;
  wire       [6:0]    _zz_when_ArraySlice_l118_283_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_283_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_283_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_283_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_283_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_283_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_283_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_283_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_283_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_283_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_284;
  wire       [5:0]    _zz_when_ArraySlice_l165_284_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_284;
  wire       [5:0]    _zz_when_ArraySlice_l166_284_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_284_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_284_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_284;
  wire       [6:0]    _zz_when_ArraySlice_l113_284;
  wire       [6:0]    _zz_when_ArraySlice_l113_284_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_284_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_284_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_284_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_284;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_284_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_284_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_284_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_284;
  wire       [6:0]    _zz_when_ArraySlice_l118_284_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_284_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_284_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_284_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_284_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_284_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_284_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_284_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_284_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_285;
  wire       [5:0]    _zz_when_ArraySlice_l165_285_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_285;
  wire       [4:0]    _zz_when_ArraySlice_l166_285_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_285_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_285_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_285_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_285;
  wire       [6:0]    _zz_when_ArraySlice_l113_285;
  wire       [6:0]    _zz_when_ArraySlice_l113_285_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_285_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_285_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_285_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_285;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_285_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_285_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_285_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_285;
  wire       [6:0]    _zz_when_ArraySlice_l118_285_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_285_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_285_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_285_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_285_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_285_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_285_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_285_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_285_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_286;
  wire       [5:0]    _zz_when_ArraySlice_l165_286_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_286;
  wire       [4:0]    _zz_when_ArraySlice_l166_286_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_286_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_286_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_286_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_286;
  wire       [6:0]    _zz_when_ArraySlice_l113_286;
  wire       [6:0]    _zz_when_ArraySlice_l113_286_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_286_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_286_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_286_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_286;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_286_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_286_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_286_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_286;
  wire       [6:0]    _zz_when_ArraySlice_l118_286_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_286_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_286_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_286_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_286_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_286_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_286_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_286_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_286_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_287;
  wire       [5:0]    _zz_when_ArraySlice_l165_287_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_287;
  wire       [3:0]    _zz_when_ArraySlice_l166_287_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_287_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_287_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_287_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_287;
  wire       [6:0]    _zz_when_ArraySlice_l113_287;
  wire       [6:0]    _zz_when_ArraySlice_l113_287_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_287_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_287_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_287_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_287;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_287_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_287_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_287_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_287;
  wire       [6:0]    _zz_when_ArraySlice_l118_287_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_287_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_287_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_287_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_287_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_287_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_287_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_287_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_287_8;
  wire                _zz_when_ArraySlice_l265_3_1;
  wire                _zz_when_ArraySlice_l265_3_2;
  wire                _zz_when_ArraySlice_l265_3_3;
  wire                _zz_when_ArraySlice_l265_3_4;
  wire                _zz_when_ArraySlice_l265_3_5;
  wire                _zz_when_ArraySlice_l265_3_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l268_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l268_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l268_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l268_3_5;
  wire       [0:0]    _zz_when_ArraySlice_l268_3_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_3_7;
  wire       [4:0]    _zz_when_ArraySlice_l268_3_8;
  wire       [5:0]    _zz_selectReadFifo_3_46;
  wire       [0:0]    _zz_selectReadFifo_3_47;
  wire       [12:0]   _zz_when_ArraySlice_l272_3_1;
  wire       [12:0]   _zz_when_ArraySlice_l272_3_2;
  wire       [12:0]   _zz_when_ArraySlice_l272_3_3;
  wire       [0:0]    _zz_when_ArraySlice_l272_3_4;
  reg        [6:0]    _zz_when_ArraySlice_l276_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l276_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l276_3_3;
  wire       [4:0]    _zz_when_ArraySlice_l276_3_4;
  wire       [12:0]   _zz_when_ArraySlice_l277_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l277_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l277_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l277_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l277_3_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_34;
  wire       [6:0]    _zz_when_ArraySlice_l95_34;
  wire       [6:0]    _zz_when_ArraySlice_l95_34_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_34_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_34_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_34_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_3_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_3_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_3_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_34;
  wire       [6:0]    _zz_when_ArraySlice_l99_34_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_3_2;
  wire       [0:0]    _zz_when_ArraySlice_l279_3_3;
  wire       [6:0]    _zz_when_ArraySlice_l279_3_4;
  wire       [5:0]    _zz_selectReadFifo_3_48;
  wire       [5:0]    _zz_selectReadFifo_3_49;
  wire       [5:0]    _zz_selectReadFifo_3_50;
  wire       [0:0]    _zz_selectReadFifo_3_51;
  wire       [5:0]    _zz_selectReadFifo_3_52;
  wire       [5:0]    _zz_selectReadFifo_3_53;
  wire       [5:0]    _zz_selectReadFifo_3_54;
  wire       [0:0]    _zz_selectReadFifo_3_55;
  wire       [5:0]    _zz_when_ArraySlice_l165_288;
  wire       [5:0]    _zz_when_ArraySlice_l165_288_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_288_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_288;
  wire       [6:0]    _zz_when_ArraySlice_l166_288_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_288_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_288_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_288_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_288_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_288;
  wire       [6:0]    _zz_when_ArraySlice_l113_288;
  wire       [6:0]    _zz_when_ArraySlice_l113_288_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_288_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_288_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_288_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_288;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_288_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_288_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_288_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_288;
  wire       [6:0]    _zz_when_ArraySlice_l118_288_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_288_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_288_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_288_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_288_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_288_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_288_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_288_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_288_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_289;
  wire       [5:0]    _zz_when_ArraySlice_l165_289_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_289_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_289;
  wire       [5:0]    _zz_when_ArraySlice_l166_289_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_289_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_289_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_289_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_289;
  wire       [6:0]    _zz_when_ArraySlice_l113_289;
  wire       [6:0]    _zz_when_ArraySlice_l113_289_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_289_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_289_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_289_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_289;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_289_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_289_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_289_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_289;
  wire       [6:0]    _zz_when_ArraySlice_l118_289_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_289_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_289_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_289_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_289_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_289_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_289_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_289_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_289_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_289_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_290;
  wire       [5:0]    _zz_when_ArraySlice_l165_290_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_290_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_290;
  wire       [5:0]    _zz_when_ArraySlice_l166_290_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_290_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_290_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_290_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_290;
  wire       [6:0]    _zz_when_ArraySlice_l113_290;
  wire       [6:0]    _zz_when_ArraySlice_l113_290_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_290_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_290_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_290_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_290;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_290_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_290_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_290_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_290;
  wire       [6:0]    _zz_when_ArraySlice_l118_290_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_290_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_290_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_290_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_290_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_290_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_290_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_290_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_290_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_290_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_291;
  wire       [5:0]    _zz_when_ArraySlice_l165_291_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_291_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_291;
  wire       [5:0]    _zz_when_ArraySlice_l166_291_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_291_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_291_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_291_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_291;
  wire       [6:0]    _zz_when_ArraySlice_l113_291;
  wire       [6:0]    _zz_when_ArraySlice_l113_291_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_291_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_291_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_291_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_291;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_291_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_291_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_291_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_291;
  wire       [6:0]    _zz_when_ArraySlice_l118_291_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_291_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_291_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_291_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_291_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_291_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_291_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_291_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_291_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_291_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_292;
  wire       [5:0]    _zz_when_ArraySlice_l165_292_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_292;
  wire       [5:0]    _zz_when_ArraySlice_l166_292_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_292_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_292_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_292;
  wire       [6:0]    _zz_when_ArraySlice_l113_292;
  wire       [6:0]    _zz_when_ArraySlice_l113_292_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_292_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_292_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_292_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_292;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_292_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_292_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_292_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_292;
  wire       [6:0]    _zz_when_ArraySlice_l118_292_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_292_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_292_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_292_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_292_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_292_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_292_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_292_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_292_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_293;
  wire       [5:0]    _zz_when_ArraySlice_l165_293_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_293;
  wire       [4:0]    _zz_when_ArraySlice_l166_293_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_293_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_293_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_293_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_293;
  wire       [6:0]    _zz_when_ArraySlice_l113_293;
  wire       [6:0]    _zz_when_ArraySlice_l113_293_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_293_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_293_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_293_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_293;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_293_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_293_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_293_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_293;
  wire       [6:0]    _zz_when_ArraySlice_l118_293_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_293_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_293_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_293_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_293_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_293_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_293_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_293_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_293_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_294;
  wire       [5:0]    _zz_when_ArraySlice_l165_294_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_294;
  wire       [4:0]    _zz_when_ArraySlice_l166_294_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_294_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_294_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_294_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_294;
  wire       [6:0]    _zz_when_ArraySlice_l113_294;
  wire       [6:0]    _zz_when_ArraySlice_l113_294_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_294_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_294_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_294_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_294;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_294_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_294_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_294_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_294;
  wire       [6:0]    _zz_when_ArraySlice_l118_294_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_294_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_294_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_294_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_294_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_294_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_294_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_294_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_294_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_295;
  wire       [5:0]    _zz_when_ArraySlice_l165_295_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_295;
  wire       [3:0]    _zz_when_ArraySlice_l166_295_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_295_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_295_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_295_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_295;
  wire       [6:0]    _zz_when_ArraySlice_l113_295;
  wire       [6:0]    _zz_when_ArraySlice_l113_295_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_295_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_295_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_295_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_295;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_295_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_295_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_295_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_295;
  wire       [6:0]    _zz_when_ArraySlice_l118_295_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_295_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_295_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_295_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_295_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_295_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_295_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_295_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_295_8;
  wire                _zz_when_ArraySlice_l285_3_1;
  wire                _zz_when_ArraySlice_l285_3_2;
  wire                _zz_when_ArraySlice_l285_3_3;
  wire                _zz_when_ArraySlice_l285_3_4;
  wire                _zz_when_ArraySlice_l285_3_5;
  wire                _zz_when_ArraySlice_l285_3_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l288_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l288_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l288_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l288_3_5;
  wire       [0:0]    _zz_when_ArraySlice_l288_3_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_3_7;
  wire       [4:0]    _zz_when_ArraySlice_l288_3_8;
  wire       [5:0]    _zz_selectReadFifo_3_56;
  wire       [0:0]    _zz_selectReadFifo_3_57;
  wire       [12:0]   _zz_when_ArraySlice_l292_3_1;
  wire       [12:0]   _zz_when_ArraySlice_l292_3_2;
  wire       [12:0]   _zz_when_ArraySlice_l292_3_3;
  wire       [0:0]    _zz_when_ArraySlice_l292_3_4;
  wire       [12:0]   _zz_when_ArraySlice_l303_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l303_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l303_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l303_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l303_3_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_35;
  wire       [6:0]    _zz_when_ArraySlice_l95_35;
  wire       [6:0]    _zz_when_ArraySlice_l95_35_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_35_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_35_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_35_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_3_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_3_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_3_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l99_35;
  wire       [6:0]    _zz_when_ArraySlice_l99_35_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_3_2;
  wire       [0:0]    _zz_when_ArraySlice_l304_3_3;
  wire       [6:0]    _zz_when_ArraySlice_l304_3_4;
  wire       [5:0]    _zz_selectReadFifo_3_58;
  wire       [5:0]    _zz_selectReadFifo_3_59;
  wire       [5:0]    _zz_selectReadFifo_3_60;
  wire       [0:0]    _zz_selectReadFifo_3_61;
  wire       [5:0]    _zz_when_ArraySlice_l165_296;
  wire       [5:0]    _zz_when_ArraySlice_l165_296_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_296_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_296;
  wire       [6:0]    _zz_when_ArraySlice_l166_296_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_296_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_296_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_296_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_296_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_296;
  wire       [6:0]    _zz_when_ArraySlice_l113_296;
  wire       [6:0]    _zz_when_ArraySlice_l113_296_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_296_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_296_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_296_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_296;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_296_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_296_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_296_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_296;
  wire       [6:0]    _zz_when_ArraySlice_l118_296_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_296_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_296_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_296_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_296_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_296_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_296_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_296_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_296_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_297;
  wire       [5:0]    _zz_when_ArraySlice_l165_297_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_297_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_297;
  wire       [5:0]    _zz_when_ArraySlice_l166_297_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_297_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_297_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_297_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_297;
  wire       [6:0]    _zz_when_ArraySlice_l113_297;
  wire       [6:0]    _zz_when_ArraySlice_l113_297_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_297_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_297_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_297_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_297;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_297_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_297_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_297_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_297;
  wire       [6:0]    _zz_when_ArraySlice_l118_297_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_297_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_297_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_297_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_297_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_297_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_297_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_297_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_297_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_297_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_298;
  wire       [5:0]    _zz_when_ArraySlice_l165_298_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_298_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_298;
  wire       [5:0]    _zz_when_ArraySlice_l166_298_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_298_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_298_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_298_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_298;
  wire       [6:0]    _zz_when_ArraySlice_l113_298;
  wire       [6:0]    _zz_when_ArraySlice_l113_298_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_298_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_298_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_298_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_298;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_298_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_298_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_298_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_298;
  wire       [6:0]    _zz_when_ArraySlice_l118_298_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_298_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_298_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_298_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_298_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_298_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_298_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_298_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_298_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_298_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_299;
  wire       [5:0]    _zz_when_ArraySlice_l165_299_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_299_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_299;
  wire       [5:0]    _zz_when_ArraySlice_l166_299_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_299_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_299_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_299_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_299;
  wire       [6:0]    _zz_when_ArraySlice_l113_299;
  wire       [6:0]    _zz_when_ArraySlice_l113_299_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_299_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_299_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_299_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_299;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_299_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_299_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_299_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_299;
  wire       [6:0]    _zz_when_ArraySlice_l118_299_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_299_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_299_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_299_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_299_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_299_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_299_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_299_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_299_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_299_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_300;
  wire       [5:0]    _zz_when_ArraySlice_l165_300_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_300;
  wire       [5:0]    _zz_when_ArraySlice_l166_300_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_300_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_300_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_300;
  wire       [6:0]    _zz_when_ArraySlice_l113_300;
  wire       [6:0]    _zz_when_ArraySlice_l113_300_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_300_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_300_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_300_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_300;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_300_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_300_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_300_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_300;
  wire       [6:0]    _zz_when_ArraySlice_l118_300_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_300_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_300_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_300_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_300_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_300_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_300_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_300_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_300_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_301;
  wire       [5:0]    _zz_when_ArraySlice_l165_301_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_301;
  wire       [4:0]    _zz_when_ArraySlice_l166_301_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_301_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_301_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_301_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_301;
  wire       [6:0]    _zz_when_ArraySlice_l113_301;
  wire       [6:0]    _zz_when_ArraySlice_l113_301_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_301_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_301_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_301_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_301;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_301_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_301_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_301_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_301;
  wire       [6:0]    _zz_when_ArraySlice_l118_301_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_301_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_301_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_301_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_301_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_301_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_301_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_301_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_301_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_302;
  wire       [5:0]    _zz_when_ArraySlice_l165_302_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_302;
  wire       [4:0]    _zz_when_ArraySlice_l166_302_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_302_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_302_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_302_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_302;
  wire       [6:0]    _zz_when_ArraySlice_l113_302;
  wire       [6:0]    _zz_when_ArraySlice_l113_302_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_302_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_302_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_302_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_302;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_302_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_302_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_302_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_302;
  wire       [6:0]    _zz_when_ArraySlice_l118_302_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_302_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_302_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_302_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_302_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_302_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_302_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_302_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_302_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_303;
  wire       [5:0]    _zz_when_ArraySlice_l165_303_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_303;
  wire       [3:0]    _zz_when_ArraySlice_l166_303_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_303_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_303_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_303_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_303;
  wire       [6:0]    _zz_when_ArraySlice_l113_303;
  wire       [6:0]    _zz_when_ArraySlice_l113_303_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_303_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_303_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_303_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_303;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_303_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_303_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_303_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_303;
  wire       [6:0]    _zz_when_ArraySlice_l118_303_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_303_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_303_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_303_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_303_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_303_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_303_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_303_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_303_8;
  wire                _zz_when_ArraySlice_l311_3_1;
  wire                _zz_when_ArraySlice_l311_3_2;
  wire                _zz_when_ArraySlice_l311_3_3;
  wire                _zz_when_ArraySlice_l311_3_4;
  wire                _zz_when_ArraySlice_l311_3_5;
  wire                _zz_when_ArraySlice_l311_3_6;
  wire       [5:0]    _zz_selectReadFifo_3_62;
  wire       [0:0]    _zz_selectReadFifo_3_63;
  wire       [12:0]   _zz_when_ArraySlice_l315_3_1;
  wire       [12:0]   _zz_when_ArraySlice_l315_3_2;
  wire       [12:0]   _zz_when_ArraySlice_l315_3_3;
  wire       [0:0]    _zz_when_ArraySlice_l315_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l301_3;
  wire       [5:0]    _zz_when_ArraySlice_l301_3_1;
  wire       [4:0]    _zz_when_ArraySlice_l301_3_2;
  wire       [12:0]   _zz_when_ArraySlice_l322_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l322_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l322_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l322_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l322_3_5;
  wire       [5:0]    _zz_when_ArraySlice_l240_4;
  wire       [5:0]    _zz_when_ArraySlice_l240_4_1;
  reg        [6:0]    _zz_when_ArraySlice_l241_4;
  wire       [5:0]    _zz_when_ArraySlice_l241_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l241_4_2;
  wire       [5:0]    _zz__zz_outputStreamArrayData_4_valid_1;
  reg                 _zz_outputStreamArrayData_4_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_4_payload_1;
  wire       [6:0]    _zz_when_ArraySlice_l247_4_1;
  wire       [0:0]    _zz_when_ArraySlice_l247_4_2;
  reg        [6:0]    _zz_when_ArraySlice_l247_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l247_4_4;
  wire       [5:0]    _zz_when_ArraySlice_l247_4_5;
  wire       [12:0]   _zz_when_ArraySlice_l248_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l248_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l248_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l248_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l248_4_5;
  wire       [5:0]    _zz_selectReadFifo_4_32;
  wire       [5:0]    _zz_selectReadFifo_4_33;
  wire       [5:0]    _zz_selectReadFifo_4_34;
  wire       [0:0]    _zz_selectReadFifo_4_35;
  wire       [5:0]    _zz_selectReadFifo_4_36;
  wire       [0:0]    _zz_selectReadFifo_4_37;
  wire       [12:0]   _zz_when_ArraySlice_l251_4;
  wire       [12:0]   _zz_when_ArraySlice_l251_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l251_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l251_4_3;
  reg        [6:0]    _zz_when_ArraySlice_l256_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l256_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l256_4_3;
  wire       [6:0]    _zz_when_ArraySlice_l256_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l256_4_5;
  wire       [12:0]   _zz_when_ArraySlice_l257_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l257_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l257_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l257_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l257_4_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_36;
  wire       [6:0]    _zz_when_ArraySlice_l95_36;
  wire       [6:0]    _zz_when_ArraySlice_l95_36_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_36_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_36_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_36_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_4_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_4_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_36;
  wire       [6:0]    _zz_when_ArraySlice_l99_36_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l259_4_3;
  wire       [6:0]    _zz_when_ArraySlice_l259_4_4;
  wire       [5:0]    _zz_selectReadFifo_4_38;
  wire       [5:0]    _zz_selectReadFifo_4_39;
  wire       [5:0]    _zz_selectReadFifo_4_40;
  wire       [0:0]    _zz_selectReadFifo_4_41;
  wire       [5:0]    _zz_selectReadFifo_4_42;
  wire       [5:0]    _zz_selectReadFifo_4_43;
  wire       [5:0]    _zz_selectReadFifo_4_44;
  wire       [0:0]    _zz_selectReadFifo_4_45;
  wire       [5:0]    _zz_when_ArraySlice_l165_304;
  wire       [5:0]    _zz_when_ArraySlice_l165_304_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_304_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_304;
  wire       [6:0]    _zz_when_ArraySlice_l166_304_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_304_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_304_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_304_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_304_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_304;
  wire       [6:0]    _zz_when_ArraySlice_l113_304;
  wire       [6:0]    _zz_when_ArraySlice_l113_304_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_304_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_304_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_304_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_304;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_304_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_304_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_304_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_304;
  wire       [6:0]    _zz_when_ArraySlice_l118_304_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_304_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_304_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_304_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_304_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_304_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_304_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_304_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_304_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_305;
  wire       [5:0]    _zz_when_ArraySlice_l165_305_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_305_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_305;
  wire       [5:0]    _zz_when_ArraySlice_l166_305_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_305_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_305_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_305_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_305;
  wire       [6:0]    _zz_when_ArraySlice_l113_305;
  wire       [6:0]    _zz_when_ArraySlice_l113_305_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_305_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_305_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_305_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_305;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_305_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_305_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_305_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_305;
  wire       [6:0]    _zz_when_ArraySlice_l118_305_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_305_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_305_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_305_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_305_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_305_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_305_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_305_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_305_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_305_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_306;
  wire       [5:0]    _zz_when_ArraySlice_l165_306_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_306_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_306;
  wire       [5:0]    _zz_when_ArraySlice_l166_306_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_306_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_306_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_306_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_306;
  wire       [6:0]    _zz_when_ArraySlice_l113_306;
  wire       [6:0]    _zz_when_ArraySlice_l113_306_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_306_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_306_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_306_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_306;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_306_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_306_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_306_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_306;
  wire       [6:0]    _zz_when_ArraySlice_l118_306_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_306_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_306_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_306_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_306_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_306_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_306_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_306_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_306_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_306_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_307;
  wire       [5:0]    _zz_when_ArraySlice_l165_307_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_307_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_307;
  wire       [5:0]    _zz_when_ArraySlice_l166_307_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_307_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_307_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_307_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_307;
  wire       [6:0]    _zz_when_ArraySlice_l113_307;
  wire       [6:0]    _zz_when_ArraySlice_l113_307_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_307_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_307_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_307_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_307;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_307_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_307_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_307_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_307;
  wire       [6:0]    _zz_when_ArraySlice_l118_307_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_307_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_307_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_307_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_307_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_307_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_307_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_307_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_307_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_307_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_308;
  wire       [5:0]    _zz_when_ArraySlice_l165_308_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_308;
  wire       [5:0]    _zz_when_ArraySlice_l166_308_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_308_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_308_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_308;
  wire       [6:0]    _zz_when_ArraySlice_l113_308;
  wire       [6:0]    _zz_when_ArraySlice_l113_308_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_308_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_308_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_308_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_308;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_308_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_308_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_308_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_308;
  wire       [6:0]    _zz_when_ArraySlice_l118_308_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_308_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_308_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_308_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_308_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_308_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_308_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_308_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_308_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_309;
  wire       [5:0]    _zz_when_ArraySlice_l165_309_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_309;
  wire       [4:0]    _zz_when_ArraySlice_l166_309_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_309_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_309_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_309_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_309;
  wire       [6:0]    _zz_when_ArraySlice_l113_309;
  wire       [6:0]    _zz_when_ArraySlice_l113_309_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_309_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_309_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_309_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_309;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_309_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_309_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_309_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_309;
  wire       [6:0]    _zz_when_ArraySlice_l118_309_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_309_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_309_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_309_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_309_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_309_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_309_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_309_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_309_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_310;
  wire       [5:0]    _zz_when_ArraySlice_l165_310_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_310;
  wire       [4:0]    _zz_when_ArraySlice_l166_310_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_310_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_310_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_310_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_310;
  wire       [6:0]    _zz_when_ArraySlice_l113_310;
  wire       [6:0]    _zz_when_ArraySlice_l113_310_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_310_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_310_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_310_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_310;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_310_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_310_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_310_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_310;
  wire       [6:0]    _zz_when_ArraySlice_l118_310_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_310_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_310_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_310_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_310_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_310_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_310_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_310_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_310_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_311;
  wire       [5:0]    _zz_when_ArraySlice_l165_311_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_311;
  wire       [3:0]    _zz_when_ArraySlice_l166_311_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_311_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_311_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_311_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_311;
  wire       [6:0]    _zz_when_ArraySlice_l113_311;
  wire       [6:0]    _zz_when_ArraySlice_l113_311_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_311_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_311_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_311_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_311;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_311_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_311_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_311_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_311;
  wire       [6:0]    _zz_when_ArraySlice_l118_311_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_311_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_311_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_311_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_311_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_311_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_311_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_311_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_311_8;
  wire                _zz_when_ArraySlice_l265_4_1;
  wire                _zz_when_ArraySlice_l265_4_2;
  wire                _zz_when_ArraySlice_l265_4_3;
  wire                _zz_when_ArraySlice_l265_4_4;
  wire                _zz_when_ArraySlice_l265_4_5;
  wire                _zz_when_ArraySlice_l265_4_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l268_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l268_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l268_4_4;
  wire       [5:0]    _zz_when_ArraySlice_l268_4_5;
  wire       [0:0]    _zz_when_ArraySlice_l268_4_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_4_7;
  wire       [5:0]    _zz_selectReadFifo_4_46;
  wire       [0:0]    _zz_selectReadFifo_4_47;
  wire       [12:0]   _zz_when_ArraySlice_l272_4;
  wire       [12:0]   _zz_when_ArraySlice_l272_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l272_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l272_4_3;
  reg        [6:0]    _zz_when_ArraySlice_l276_4;
  wire       [5:0]    _zz_when_ArraySlice_l276_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l276_4_2;
  wire       [12:0]   _zz_when_ArraySlice_l277_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l277_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l277_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l277_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l277_4_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_37;
  wire       [6:0]    _zz_when_ArraySlice_l95_37;
  wire       [6:0]    _zz_when_ArraySlice_l95_37_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_37_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_37_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_37_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_4_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_4_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_37;
  wire       [6:0]    _zz_when_ArraySlice_l99_37_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l279_4_3;
  wire       [6:0]    _zz_when_ArraySlice_l279_4_4;
  wire       [5:0]    _zz_selectReadFifo_4_48;
  wire       [5:0]    _zz_selectReadFifo_4_49;
  wire       [5:0]    _zz_selectReadFifo_4_50;
  wire       [0:0]    _zz_selectReadFifo_4_51;
  wire       [5:0]    _zz_selectReadFifo_4_52;
  wire       [5:0]    _zz_selectReadFifo_4_53;
  wire       [5:0]    _zz_selectReadFifo_4_54;
  wire       [0:0]    _zz_selectReadFifo_4_55;
  wire       [5:0]    _zz_when_ArraySlice_l165_312;
  wire       [5:0]    _zz_when_ArraySlice_l165_312_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_312_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_312;
  wire       [6:0]    _zz_when_ArraySlice_l166_312_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_312_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_312_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_312_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_312_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_312;
  wire       [6:0]    _zz_when_ArraySlice_l113_312;
  wire       [6:0]    _zz_when_ArraySlice_l113_312_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_312_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_312_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_312_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_312;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_312_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_312_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_312_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_312;
  wire       [6:0]    _zz_when_ArraySlice_l118_312_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_312_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_312_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_312_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_312_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_312_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_312_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_312_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_312_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_313;
  wire       [5:0]    _zz_when_ArraySlice_l165_313_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_313_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_313;
  wire       [5:0]    _zz_when_ArraySlice_l166_313_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_313_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_313_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_313_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_313;
  wire       [6:0]    _zz_when_ArraySlice_l113_313;
  wire       [6:0]    _zz_when_ArraySlice_l113_313_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_313_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_313_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_313_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_313;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_313_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_313_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_313_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_313;
  wire       [6:0]    _zz_when_ArraySlice_l118_313_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_313_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_313_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_313_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_313_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_313_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_313_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_313_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_313_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_313_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_314;
  wire       [5:0]    _zz_when_ArraySlice_l165_314_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_314_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_314;
  wire       [5:0]    _zz_when_ArraySlice_l166_314_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_314_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_314_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_314_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_314;
  wire       [6:0]    _zz_when_ArraySlice_l113_314;
  wire       [6:0]    _zz_when_ArraySlice_l113_314_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_314_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_314_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_314_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_314;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_314_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_314_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_314_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_314;
  wire       [6:0]    _zz_when_ArraySlice_l118_314_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_314_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_314_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_314_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_314_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_314_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_314_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_314_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_314_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_314_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_315;
  wire       [5:0]    _zz_when_ArraySlice_l165_315_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_315_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_315;
  wire       [5:0]    _zz_when_ArraySlice_l166_315_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_315_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_315_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_315_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_315;
  wire       [6:0]    _zz_when_ArraySlice_l113_315;
  wire       [6:0]    _zz_when_ArraySlice_l113_315_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_315_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_315_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_315_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_315;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_315_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_315_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_315_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_315;
  wire       [6:0]    _zz_when_ArraySlice_l118_315_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_315_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_315_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_315_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_315_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_315_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_315_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_315_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_315_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_315_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_316;
  wire       [5:0]    _zz_when_ArraySlice_l165_316_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_316;
  wire       [5:0]    _zz_when_ArraySlice_l166_316_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_316_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_316_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_316;
  wire       [6:0]    _zz_when_ArraySlice_l113_316;
  wire       [6:0]    _zz_when_ArraySlice_l113_316_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_316_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_316_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_316_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_316;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_316_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_316_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_316_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_316;
  wire       [6:0]    _zz_when_ArraySlice_l118_316_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_316_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_316_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_316_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_316_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_316_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_316_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_316_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_316_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_317;
  wire       [5:0]    _zz_when_ArraySlice_l165_317_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_317;
  wire       [4:0]    _zz_when_ArraySlice_l166_317_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_317_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_317_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_317_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_317;
  wire       [6:0]    _zz_when_ArraySlice_l113_317;
  wire       [6:0]    _zz_when_ArraySlice_l113_317_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_317_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_317_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_317_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_317;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_317_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_317_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_317_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_317;
  wire       [6:0]    _zz_when_ArraySlice_l118_317_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_317_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_317_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_317_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_317_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_317_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_317_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_317_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_317_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_318;
  wire       [5:0]    _zz_when_ArraySlice_l165_318_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_318;
  wire       [4:0]    _zz_when_ArraySlice_l166_318_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_318_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_318_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_318_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_318;
  wire       [6:0]    _zz_when_ArraySlice_l113_318;
  wire       [6:0]    _zz_when_ArraySlice_l113_318_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_318_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_318_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_318_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_318;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_318_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_318_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_318_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_318;
  wire       [6:0]    _zz_when_ArraySlice_l118_318_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_318_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_318_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_318_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_318_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_318_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_318_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_318_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_318_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_319;
  wire       [5:0]    _zz_when_ArraySlice_l165_319_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_319;
  wire       [3:0]    _zz_when_ArraySlice_l166_319_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_319_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_319_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_319_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_319;
  wire       [6:0]    _zz_when_ArraySlice_l113_319;
  wire       [6:0]    _zz_when_ArraySlice_l113_319_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_319_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_319_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_319_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_319;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_319_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_319_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_319_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_319;
  wire       [6:0]    _zz_when_ArraySlice_l118_319_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_319_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_319_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_319_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_319_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_319_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_319_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_319_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_319_8;
  wire                _zz_when_ArraySlice_l285_4_1;
  wire                _zz_when_ArraySlice_l285_4_2;
  wire                _zz_when_ArraySlice_l285_4_3;
  wire                _zz_when_ArraySlice_l285_4_4;
  wire                _zz_when_ArraySlice_l285_4_5;
  wire                _zz_when_ArraySlice_l285_4_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l288_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l288_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l288_4_4;
  wire       [5:0]    _zz_when_ArraySlice_l288_4_5;
  wire       [0:0]    _zz_when_ArraySlice_l288_4_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_4_7;
  wire       [5:0]    _zz_selectReadFifo_4_56;
  wire       [0:0]    _zz_selectReadFifo_4_57;
  wire       [12:0]   _zz_when_ArraySlice_l292_4;
  wire       [12:0]   _zz_when_ArraySlice_l292_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l292_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l292_4_3;
  wire       [12:0]   _zz_when_ArraySlice_l303_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l303_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l303_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l303_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l303_4_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_38;
  wire       [6:0]    _zz_when_ArraySlice_l95_38;
  wire       [6:0]    _zz_when_ArraySlice_l95_38_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_38_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_38_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_38_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_4_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_4_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_38;
  wire       [6:0]    _zz_when_ArraySlice_l99_38_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l304_4_3;
  wire       [6:0]    _zz_when_ArraySlice_l304_4_4;
  wire       [5:0]    _zz_selectReadFifo_4_58;
  wire       [5:0]    _zz_selectReadFifo_4_59;
  wire       [5:0]    _zz_selectReadFifo_4_60;
  wire       [0:0]    _zz_selectReadFifo_4_61;
  wire       [5:0]    _zz_when_ArraySlice_l165_320;
  wire       [5:0]    _zz_when_ArraySlice_l165_320_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_320_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_320;
  wire       [6:0]    _zz_when_ArraySlice_l166_320_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_320_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_320_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_320_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_320_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_320;
  wire       [6:0]    _zz_when_ArraySlice_l113_320;
  wire       [6:0]    _zz_when_ArraySlice_l113_320_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_320_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_320_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_320_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_320;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_320_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_320_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_320_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_320;
  wire       [6:0]    _zz_when_ArraySlice_l118_320_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_320_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_320_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_320_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_320_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_320_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_320_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_320_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_320_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_321;
  wire       [5:0]    _zz_when_ArraySlice_l165_321_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_321_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_321;
  wire       [5:0]    _zz_when_ArraySlice_l166_321_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_321_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_321_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_321_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_321;
  wire       [6:0]    _zz_when_ArraySlice_l113_321;
  wire       [6:0]    _zz_when_ArraySlice_l113_321_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_321_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_321_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_321_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_321;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_321_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_321_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_321_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_321;
  wire       [6:0]    _zz_when_ArraySlice_l118_321_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_321_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_321_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_321_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_321_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_321_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_321_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_321_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_321_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_321_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_322;
  wire       [5:0]    _zz_when_ArraySlice_l165_322_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_322_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_322;
  wire       [5:0]    _zz_when_ArraySlice_l166_322_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_322_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_322_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_322_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_322;
  wire       [6:0]    _zz_when_ArraySlice_l113_322;
  wire       [6:0]    _zz_when_ArraySlice_l113_322_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_322_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_322_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_322_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_322;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_322_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_322_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_322_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_322;
  wire       [6:0]    _zz_when_ArraySlice_l118_322_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_322_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_322_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_322_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_322_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_322_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_322_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_322_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_322_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_322_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_323;
  wire       [5:0]    _zz_when_ArraySlice_l165_323_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_323_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_323;
  wire       [5:0]    _zz_when_ArraySlice_l166_323_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_323_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_323_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_323_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_323;
  wire       [6:0]    _zz_when_ArraySlice_l113_323;
  wire       [6:0]    _zz_when_ArraySlice_l113_323_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_323_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_323_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_323_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_323;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_323_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_323_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_323_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_323;
  wire       [6:0]    _zz_when_ArraySlice_l118_323_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_323_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_323_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_323_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_323_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_323_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_323_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_323_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_323_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_323_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_324;
  wire       [5:0]    _zz_when_ArraySlice_l165_324_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_324;
  wire       [5:0]    _zz_when_ArraySlice_l166_324_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_324_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_324_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_324;
  wire       [6:0]    _zz_when_ArraySlice_l113_324;
  wire       [6:0]    _zz_when_ArraySlice_l113_324_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_324_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_324_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_324_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_324;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_324_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_324_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_324_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_324;
  wire       [6:0]    _zz_when_ArraySlice_l118_324_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_324_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_324_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_324_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_324_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_324_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_324_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_324_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_324_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_325;
  wire       [5:0]    _zz_when_ArraySlice_l165_325_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_325;
  wire       [4:0]    _zz_when_ArraySlice_l166_325_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_325_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_325_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_325_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_325;
  wire       [6:0]    _zz_when_ArraySlice_l113_325;
  wire       [6:0]    _zz_when_ArraySlice_l113_325_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_325_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_325_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_325_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_325;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_325_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_325_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_325_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_325;
  wire       [6:0]    _zz_when_ArraySlice_l118_325_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_325_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_325_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_325_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_325_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_325_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_325_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_325_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_325_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_326;
  wire       [5:0]    _zz_when_ArraySlice_l165_326_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_326;
  wire       [4:0]    _zz_when_ArraySlice_l166_326_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_326_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_326_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_326_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_326;
  wire       [6:0]    _zz_when_ArraySlice_l113_326;
  wire       [6:0]    _zz_when_ArraySlice_l113_326_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_326_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_326_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_326_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_326;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_326_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_326_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_326_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_326;
  wire       [6:0]    _zz_when_ArraySlice_l118_326_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_326_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_326_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_326_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_326_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_326_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_326_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_326_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_326_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_327;
  wire       [5:0]    _zz_when_ArraySlice_l165_327_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_327;
  wire       [3:0]    _zz_when_ArraySlice_l166_327_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_327_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_327_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_327_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_327;
  wire       [6:0]    _zz_when_ArraySlice_l113_327;
  wire       [6:0]    _zz_when_ArraySlice_l113_327_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_327_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_327_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_327_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_327;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_327_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_327_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_327_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_327;
  wire       [6:0]    _zz_when_ArraySlice_l118_327_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_327_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_327_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_327_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_327_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_327_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_327_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_327_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_327_8;
  wire                _zz_when_ArraySlice_l311_4_1;
  wire                _zz_when_ArraySlice_l311_4_2;
  wire                _zz_when_ArraySlice_l311_4_3;
  wire                _zz_when_ArraySlice_l311_4_4;
  wire                _zz_when_ArraySlice_l311_4_5;
  wire                _zz_when_ArraySlice_l311_4_6;
  wire       [5:0]    _zz_selectReadFifo_4_62;
  wire       [0:0]    _zz_selectReadFifo_4_63;
  wire       [12:0]   _zz_when_ArraySlice_l315_4;
  wire       [12:0]   _zz_when_ArraySlice_l315_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l315_4_2;
  wire       [0:0]    _zz_when_ArraySlice_l315_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l301_4;
  wire       [5:0]    _zz_when_ArraySlice_l301_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l322_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l322_4_2;
  wire       [5:0]    _zz_when_ArraySlice_l322_4_3;
  wire       [5:0]    _zz_when_ArraySlice_l322_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l322_4_5;
  wire       [5:0]    _zz_when_ArraySlice_l240_5;
  wire       [5:0]    _zz_when_ArraySlice_l240_5_1;
  reg        [6:0]    _zz_when_ArraySlice_l241_5;
  wire       [5:0]    _zz_when_ArraySlice_l241_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l241_5_2;
  wire       [5:0]    _zz__zz_outputStreamArrayData_5_valid_1;
  reg                 _zz_outputStreamArrayData_5_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_5_payload_1;
  wire       [6:0]    _zz_when_ArraySlice_l247_5_1;
  wire       [0:0]    _zz_when_ArraySlice_l247_5_2;
  reg        [6:0]    _zz_when_ArraySlice_l247_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l247_5_4;
  wire       [5:0]    _zz_when_ArraySlice_l247_5_5;
  wire       [12:0]   _zz_when_ArraySlice_l248_5;
  wire       [5:0]    _zz_when_ArraySlice_l248_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l248_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l248_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l248_5_4;
  wire       [5:0]    _zz_selectReadFifo_5_32;
  wire       [5:0]    _zz_selectReadFifo_5_33;
  wire       [5:0]    _zz_selectReadFifo_5_34;
  wire       [0:0]    _zz_selectReadFifo_5_35;
  wire       [5:0]    _zz_selectReadFifo_5_36;
  wire       [0:0]    _zz_selectReadFifo_5_37;
  wire       [12:0]   _zz_when_ArraySlice_l251_5;
  wire       [12:0]   _zz_when_ArraySlice_l251_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l251_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l251_5_3;
  reg        [6:0]    _zz_when_ArraySlice_l256_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l256_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l256_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l256_5_4;
  wire       [0:0]    _zz_when_ArraySlice_l256_5_5;
  wire       [12:0]   _zz_when_ArraySlice_l257_5;
  wire       [5:0]    _zz_when_ArraySlice_l257_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l257_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l257_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l257_5_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_39;
  wire       [6:0]    _zz_when_ArraySlice_l95_39;
  wire       [6:0]    _zz_when_ArraySlice_l95_39_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_39_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_39_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_39_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_5_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_5_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_39;
  wire       [6:0]    _zz_when_ArraySlice_l99_39_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l259_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l259_5_4;
  wire       [5:0]    _zz_selectReadFifo_5_38;
  wire       [5:0]    _zz_selectReadFifo_5_39;
  wire       [5:0]    _zz_selectReadFifo_5_40;
  wire       [0:0]    _zz_selectReadFifo_5_41;
  wire       [5:0]    _zz_selectReadFifo_5_42;
  wire       [5:0]    _zz_selectReadFifo_5_43;
  wire       [5:0]    _zz_selectReadFifo_5_44;
  wire       [0:0]    _zz_selectReadFifo_5_45;
  wire       [5:0]    _zz_when_ArraySlice_l165_328;
  wire       [5:0]    _zz_when_ArraySlice_l165_328_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_328_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_328;
  wire       [6:0]    _zz_when_ArraySlice_l166_328_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_328_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_328_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_328_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_328_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_328;
  wire       [6:0]    _zz_when_ArraySlice_l113_328;
  wire       [6:0]    _zz_when_ArraySlice_l113_328_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_328_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_328_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_328_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_328;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_328_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_328_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_328_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_328;
  wire       [6:0]    _zz_when_ArraySlice_l118_328_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_328_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_328_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_328_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_328_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_328_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_328_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_328_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_328_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_329;
  wire       [5:0]    _zz_when_ArraySlice_l165_329_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_329_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_329;
  wire       [5:0]    _zz_when_ArraySlice_l166_329_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_329_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_329_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_329_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_329;
  wire       [6:0]    _zz_when_ArraySlice_l113_329;
  wire       [6:0]    _zz_when_ArraySlice_l113_329_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_329_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_329_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_329_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_329;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_329_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_329_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_329_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_329;
  wire       [6:0]    _zz_when_ArraySlice_l118_329_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_329_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_329_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_329_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_329_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_329_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_329_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_329_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_329_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_329_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_330;
  wire       [5:0]    _zz_when_ArraySlice_l165_330_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_330_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_330;
  wire       [5:0]    _zz_when_ArraySlice_l166_330_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_330_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_330_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_330_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_330;
  wire       [6:0]    _zz_when_ArraySlice_l113_330;
  wire       [6:0]    _zz_when_ArraySlice_l113_330_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_330_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_330_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_330_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_330;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_330_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_330_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_330_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_330;
  wire       [6:0]    _zz_when_ArraySlice_l118_330_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_330_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_330_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_330_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_330_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_330_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_330_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_330_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_330_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_330_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_331;
  wire       [5:0]    _zz_when_ArraySlice_l165_331_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_331_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_331;
  wire       [5:0]    _zz_when_ArraySlice_l166_331_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_331_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_331_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_331_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_331;
  wire       [6:0]    _zz_when_ArraySlice_l113_331;
  wire       [6:0]    _zz_when_ArraySlice_l113_331_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_331_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_331_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_331_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_331;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_331_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_331_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_331_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_331;
  wire       [6:0]    _zz_when_ArraySlice_l118_331_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_331_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_331_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_331_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_331_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_331_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_331_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_331_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_331_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_331_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_332;
  wire       [5:0]    _zz_when_ArraySlice_l165_332_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_332;
  wire       [5:0]    _zz_when_ArraySlice_l166_332_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_332_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_332_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_332;
  wire       [6:0]    _zz_when_ArraySlice_l113_332;
  wire       [6:0]    _zz_when_ArraySlice_l113_332_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_332_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_332_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_332_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_332;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_332_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_332_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_332_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_332;
  wire       [6:0]    _zz_when_ArraySlice_l118_332_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_332_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_332_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_332_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_332_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_332_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_332_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_332_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_332_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_333;
  wire       [5:0]    _zz_when_ArraySlice_l165_333_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_333;
  wire       [4:0]    _zz_when_ArraySlice_l166_333_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_333_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_333_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_333_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_333;
  wire       [6:0]    _zz_when_ArraySlice_l113_333;
  wire       [6:0]    _zz_when_ArraySlice_l113_333_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_333_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_333_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_333_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_333;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_333_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_333_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_333_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_333;
  wire       [6:0]    _zz_when_ArraySlice_l118_333_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_333_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_333_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_333_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_333_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_333_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_333_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_333_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_333_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_334;
  wire       [5:0]    _zz_when_ArraySlice_l165_334_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_334;
  wire       [4:0]    _zz_when_ArraySlice_l166_334_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_334_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_334_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_334_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_334;
  wire       [6:0]    _zz_when_ArraySlice_l113_334;
  wire       [6:0]    _zz_when_ArraySlice_l113_334_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_334_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_334_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_334_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_334;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_334_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_334_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_334_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_334;
  wire       [6:0]    _zz_when_ArraySlice_l118_334_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_334_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_334_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_334_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_334_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_334_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_334_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_334_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_334_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_335;
  wire       [5:0]    _zz_when_ArraySlice_l165_335_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_335;
  wire       [3:0]    _zz_when_ArraySlice_l166_335_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_335_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_335_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_335_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_335;
  wire       [6:0]    _zz_when_ArraySlice_l113_335;
  wire       [6:0]    _zz_when_ArraySlice_l113_335_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_335_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_335_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_335_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_335;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_335_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_335_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_335_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_335;
  wire       [6:0]    _zz_when_ArraySlice_l118_335_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_335_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_335_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_335_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_335_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_335_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_335_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_335_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_335_8;
  wire                _zz_when_ArraySlice_l265_5_1;
  wire                _zz_when_ArraySlice_l265_5_2;
  wire                _zz_when_ArraySlice_l265_5_3;
  wire                _zz_when_ArraySlice_l265_5_4;
  wire                _zz_when_ArraySlice_l265_5_5;
  wire                _zz_when_ArraySlice_l265_5_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l268_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l268_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l268_5_4;
  wire       [5:0]    _zz_when_ArraySlice_l268_5_5;
  wire       [0:0]    _zz_when_ArraySlice_l268_5_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_5_7;
  wire       [5:0]    _zz_selectReadFifo_5_46;
  wire       [0:0]    _zz_selectReadFifo_5_47;
  wire       [12:0]   _zz_when_ArraySlice_l272_5;
  wire       [12:0]   _zz_when_ArraySlice_l272_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l272_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l272_5_3;
  reg        [6:0]    _zz_when_ArraySlice_l276_5;
  wire       [5:0]    _zz_when_ArraySlice_l276_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l276_5_2;
  wire       [12:0]   _zz_when_ArraySlice_l277_5;
  wire       [5:0]    _zz_when_ArraySlice_l277_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l277_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l277_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l277_5_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_40;
  wire       [6:0]    _zz_when_ArraySlice_l95_40;
  wire       [6:0]    _zz_when_ArraySlice_l95_40_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_40_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_40_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_40_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_5_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_5_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_40;
  wire       [6:0]    _zz_when_ArraySlice_l99_40_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l279_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l279_5_4;
  wire       [5:0]    _zz_selectReadFifo_5_48;
  wire       [5:0]    _zz_selectReadFifo_5_49;
  wire       [5:0]    _zz_selectReadFifo_5_50;
  wire       [0:0]    _zz_selectReadFifo_5_51;
  wire       [5:0]    _zz_selectReadFifo_5_52;
  wire       [5:0]    _zz_selectReadFifo_5_53;
  wire       [5:0]    _zz_selectReadFifo_5_54;
  wire       [0:0]    _zz_selectReadFifo_5_55;
  wire       [5:0]    _zz_when_ArraySlice_l165_336;
  wire       [5:0]    _zz_when_ArraySlice_l165_336_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_336_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_336;
  wire       [6:0]    _zz_when_ArraySlice_l166_336_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_336_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_336_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_336_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_336_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_336;
  wire       [6:0]    _zz_when_ArraySlice_l113_336;
  wire       [6:0]    _zz_when_ArraySlice_l113_336_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_336_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_336_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_336_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_336;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_336_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_336_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_336_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_336;
  wire       [6:0]    _zz_when_ArraySlice_l118_336_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_336_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_336_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_336_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_336_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_336_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_336_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_336_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_336_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_337;
  wire       [5:0]    _zz_when_ArraySlice_l165_337_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_337_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_337;
  wire       [5:0]    _zz_when_ArraySlice_l166_337_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_337_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_337_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_337_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_337;
  wire       [6:0]    _zz_when_ArraySlice_l113_337;
  wire       [6:0]    _zz_when_ArraySlice_l113_337_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_337_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_337_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_337_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_337;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_337_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_337_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_337_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_337;
  wire       [6:0]    _zz_when_ArraySlice_l118_337_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_337_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_337_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_337_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_337_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_337_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_337_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_337_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_337_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_337_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_338;
  wire       [5:0]    _zz_when_ArraySlice_l165_338_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_338_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_338;
  wire       [5:0]    _zz_when_ArraySlice_l166_338_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_338_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_338_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_338_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_338;
  wire       [6:0]    _zz_when_ArraySlice_l113_338;
  wire       [6:0]    _zz_when_ArraySlice_l113_338_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_338_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_338_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_338_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_338;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_338_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_338_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_338_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_338;
  wire       [6:0]    _zz_when_ArraySlice_l118_338_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_338_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_338_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_338_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_338_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_338_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_338_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_338_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_338_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_338_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_339;
  wire       [5:0]    _zz_when_ArraySlice_l165_339_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_339_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_339;
  wire       [5:0]    _zz_when_ArraySlice_l166_339_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_339_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_339_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_339_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_339;
  wire       [6:0]    _zz_when_ArraySlice_l113_339;
  wire       [6:0]    _zz_when_ArraySlice_l113_339_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_339_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_339_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_339_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_339;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_339_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_339_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_339_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_339;
  wire       [6:0]    _zz_when_ArraySlice_l118_339_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_339_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_339_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_339_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_339_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_339_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_339_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_339_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_339_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_339_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_340;
  wire       [5:0]    _zz_when_ArraySlice_l165_340_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_340;
  wire       [5:0]    _zz_when_ArraySlice_l166_340_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_340_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_340_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_340;
  wire       [6:0]    _zz_when_ArraySlice_l113_340;
  wire       [6:0]    _zz_when_ArraySlice_l113_340_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_340_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_340_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_340_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_340;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_340_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_340_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_340_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_340;
  wire       [6:0]    _zz_when_ArraySlice_l118_340_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_340_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_340_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_340_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_340_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_340_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_340_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_340_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_340_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_341;
  wire       [5:0]    _zz_when_ArraySlice_l165_341_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_341;
  wire       [4:0]    _zz_when_ArraySlice_l166_341_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_341_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_341_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_341_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_341;
  wire       [6:0]    _zz_when_ArraySlice_l113_341;
  wire       [6:0]    _zz_when_ArraySlice_l113_341_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_341_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_341_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_341_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_341;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_341_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_341_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_341_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_341;
  wire       [6:0]    _zz_when_ArraySlice_l118_341_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_341_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_341_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_341_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_341_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_341_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_341_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_341_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_341_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_342;
  wire       [5:0]    _zz_when_ArraySlice_l165_342_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_342;
  wire       [4:0]    _zz_when_ArraySlice_l166_342_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_342_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_342_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_342_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_342;
  wire       [6:0]    _zz_when_ArraySlice_l113_342;
  wire       [6:0]    _zz_when_ArraySlice_l113_342_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_342_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_342_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_342_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_342;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_342_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_342_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_342_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_342;
  wire       [6:0]    _zz_when_ArraySlice_l118_342_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_342_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_342_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_342_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_342_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_342_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_342_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_342_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_342_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_343;
  wire       [5:0]    _zz_when_ArraySlice_l165_343_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_343;
  wire       [3:0]    _zz_when_ArraySlice_l166_343_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_343_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_343_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_343_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_343;
  wire       [6:0]    _zz_when_ArraySlice_l113_343;
  wire       [6:0]    _zz_when_ArraySlice_l113_343_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_343_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_343_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_343_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_343;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_343_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_343_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_343_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_343;
  wire       [6:0]    _zz_when_ArraySlice_l118_343_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_343_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_343_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_343_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_343_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_343_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_343_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_343_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_343_8;
  wire                _zz_when_ArraySlice_l285_5_1;
  wire                _zz_when_ArraySlice_l285_5_2;
  wire                _zz_when_ArraySlice_l285_5_3;
  wire                _zz_when_ArraySlice_l285_5_4;
  wire                _zz_when_ArraySlice_l285_5_5;
  wire                _zz_when_ArraySlice_l285_5_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l288_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l288_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l288_5_4;
  wire       [5:0]    _zz_when_ArraySlice_l288_5_5;
  wire       [0:0]    _zz_when_ArraySlice_l288_5_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_5_7;
  wire       [5:0]    _zz_selectReadFifo_5_56;
  wire       [0:0]    _zz_selectReadFifo_5_57;
  wire       [12:0]   _zz_when_ArraySlice_l292_5;
  wire       [12:0]   _zz_when_ArraySlice_l292_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l292_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l292_5_3;
  wire       [12:0]   _zz_when_ArraySlice_l303_5;
  wire       [5:0]    _zz_when_ArraySlice_l303_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l303_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l303_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l303_5_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_41;
  wire       [6:0]    _zz_when_ArraySlice_l95_41;
  wire       [6:0]    _zz_when_ArraySlice_l95_41_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_41_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_41_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_41_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_5_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_5_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_41;
  wire       [6:0]    _zz_when_ArraySlice_l99_41_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l304_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l304_5_4;
  wire       [5:0]    _zz_selectReadFifo_5_58;
  wire       [5:0]    _zz_selectReadFifo_5_59;
  wire       [5:0]    _zz_selectReadFifo_5_60;
  wire       [0:0]    _zz_selectReadFifo_5_61;
  wire       [5:0]    _zz_when_ArraySlice_l165_344;
  wire       [5:0]    _zz_when_ArraySlice_l165_344_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_344_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_344;
  wire       [6:0]    _zz_when_ArraySlice_l166_344_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_344_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_344_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_344_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_344_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_344;
  wire       [6:0]    _zz_when_ArraySlice_l113_344;
  wire       [6:0]    _zz_when_ArraySlice_l113_344_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_344_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_344_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_344_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_344;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_344_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_344_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_344_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_344;
  wire       [6:0]    _zz_when_ArraySlice_l118_344_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_344_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_344_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_344_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_344_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_344_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_344_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_344_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_344_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_345;
  wire       [5:0]    _zz_when_ArraySlice_l165_345_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_345_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_345;
  wire       [5:0]    _zz_when_ArraySlice_l166_345_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_345_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_345_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_345_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_345;
  wire       [6:0]    _zz_when_ArraySlice_l113_345;
  wire       [6:0]    _zz_when_ArraySlice_l113_345_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_345_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_345_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_345_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_345;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_345_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_345_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_345_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_345;
  wire       [6:0]    _zz_when_ArraySlice_l118_345_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_345_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_345_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_345_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_345_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_345_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_345_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_345_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_345_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_345_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_346;
  wire       [5:0]    _zz_when_ArraySlice_l165_346_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_346_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_346;
  wire       [5:0]    _zz_when_ArraySlice_l166_346_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_346_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_346_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_346_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_346;
  wire       [6:0]    _zz_when_ArraySlice_l113_346;
  wire       [6:0]    _zz_when_ArraySlice_l113_346_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_346_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_346_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_346_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_346;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_346_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_346_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_346_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_346;
  wire       [6:0]    _zz_when_ArraySlice_l118_346_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_346_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_346_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_346_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_346_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_346_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_346_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_346_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_346_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_346_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_347;
  wire       [5:0]    _zz_when_ArraySlice_l165_347_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_347_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_347;
  wire       [5:0]    _zz_when_ArraySlice_l166_347_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_347_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_347_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_347_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_347;
  wire       [6:0]    _zz_when_ArraySlice_l113_347;
  wire       [6:0]    _zz_when_ArraySlice_l113_347_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_347_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_347_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_347_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_347;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_347_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_347_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_347_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_347;
  wire       [6:0]    _zz_when_ArraySlice_l118_347_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_347_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_347_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_347_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_347_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_347_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_347_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_347_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_347_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_347_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_348;
  wire       [5:0]    _zz_when_ArraySlice_l165_348_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_348;
  wire       [5:0]    _zz_when_ArraySlice_l166_348_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_348_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_348_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_348;
  wire       [6:0]    _zz_when_ArraySlice_l113_348;
  wire       [6:0]    _zz_when_ArraySlice_l113_348_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_348_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_348_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_348_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_348;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_348_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_348_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_348_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_348;
  wire       [6:0]    _zz_when_ArraySlice_l118_348_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_348_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_348_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_348_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_348_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_348_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_348_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_348_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_348_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_349;
  wire       [5:0]    _zz_when_ArraySlice_l165_349_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_349;
  wire       [4:0]    _zz_when_ArraySlice_l166_349_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_349_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_349_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_349_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_349;
  wire       [6:0]    _zz_when_ArraySlice_l113_349;
  wire       [6:0]    _zz_when_ArraySlice_l113_349_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_349_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_349_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_349_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_349;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_349_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_349_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_349_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_349;
  wire       [6:0]    _zz_when_ArraySlice_l118_349_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_349_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_349_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_349_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_349_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_349_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_349_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_349_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_349_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_350;
  wire       [5:0]    _zz_when_ArraySlice_l165_350_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_350;
  wire       [4:0]    _zz_when_ArraySlice_l166_350_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_350_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_350_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_350_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_350;
  wire       [6:0]    _zz_when_ArraySlice_l113_350;
  wire       [6:0]    _zz_when_ArraySlice_l113_350_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_350_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_350_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_350_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_350;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_350_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_350_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_350_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_350;
  wire       [6:0]    _zz_when_ArraySlice_l118_350_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_350_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_350_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_350_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_350_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_350_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_350_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_350_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_350_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_351;
  wire       [5:0]    _zz_when_ArraySlice_l165_351_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_351;
  wire       [3:0]    _zz_when_ArraySlice_l166_351_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_351_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_351_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_351_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_351;
  wire       [6:0]    _zz_when_ArraySlice_l113_351;
  wire       [6:0]    _zz_when_ArraySlice_l113_351_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_351_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_351_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_351_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_351;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_351_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_351_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_351_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_351;
  wire       [6:0]    _zz_when_ArraySlice_l118_351_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_351_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_351_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_351_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_351_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_351_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_351_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_351_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_351_8;
  wire                _zz_when_ArraySlice_l311_5_1;
  wire                _zz_when_ArraySlice_l311_5_2;
  wire                _zz_when_ArraySlice_l311_5_3;
  wire                _zz_when_ArraySlice_l311_5_4;
  wire                _zz_when_ArraySlice_l311_5_5;
  wire                _zz_when_ArraySlice_l311_5_6;
  wire       [5:0]    _zz_selectReadFifo_5_62;
  wire       [0:0]    _zz_selectReadFifo_5_63;
  wire       [12:0]   _zz_when_ArraySlice_l315_5;
  wire       [12:0]   _zz_when_ArraySlice_l315_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l315_5_2;
  wire       [0:0]    _zz_when_ArraySlice_l315_5_3;
  wire       [5:0]    _zz_when_ArraySlice_l301_5;
  wire       [5:0]    _zz_when_ArraySlice_l301_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l322_5;
  wire       [5:0]    _zz_when_ArraySlice_l322_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l322_5_2;
  wire       [5:0]    _zz_when_ArraySlice_l322_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l322_5_4;
  wire       [5:0]    _zz_when_ArraySlice_l240_6;
  wire       [5:0]    _zz_when_ArraySlice_l240_6_1;
  reg        [6:0]    _zz_when_ArraySlice_l241_6;
  wire       [5:0]    _zz_when_ArraySlice_l241_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l241_6_2;
  wire       [5:0]    _zz__zz_outputStreamArrayData_6_valid_1;
  reg                 _zz_outputStreamArrayData_6_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_6_payload_1;
  wire       [6:0]    _zz_when_ArraySlice_l247_6;
  wire       [0:0]    _zz_when_ArraySlice_l247_6_1;
  reg        [6:0]    _zz_when_ArraySlice_l247_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l247_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l247_6_4;
  wire       [12:0]   _zz_when_ArraySlice_l248_6;
  wire       [5:0]    _zz_when_ArraySlice_l248_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l248_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l248_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l248_6_4;
  wire       [5:0]    _zz_selectReadFifo_6_32;
  wire       [5:0]    _zz_selectReadFifo_6_33;
  wire       [5:0]    _zz_selectReadFifo_6_34;
  wire       [0:0]    _zz_selectReadFifo_6_35;
  wire       [5:0]    _zz_selectReadFifo_6_36;
  wire       [0:0]    _zz_selectReadFifo_6_37;
  wire       [12:0]   _zz_when_ArraySlice_l251_6;
  wire       [12:0]   _zz_when_ArraySlice_l251_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l251_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l251_6_3;
  reg        [6:0]    _zz_when_ArraySlice_l256_6;
  wire       [5:0]    _zz_when_ArraySlice_l256_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l256_6_2;
  wire       [6:0]    _zz_when_ArraySlice_l256_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l256_6_4;
  wire       [12:0]   _zz_when_ArraySlice_l257_6;
  wire       [5:0]    _zz_when_ArraySlice_l257_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l257_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l257_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l257_6_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_42;
  wire       [6:0]    _zz_when_ArraySlice_l95_42;
  wire       [6:0]    _zz_when_ArraySlice_l95_42_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_42_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_42_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_42_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_6;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_6_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_6_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_42;
  wire       [6:0]    _zz_when_ArraySlice_l99_42_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l259_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l259_6_4;
  wire       [5:0]    _zz_selectReadFifo_6_38;
  wire       [5:0]    _zz_selectReadFifo_6_39;
  wire       [5:0]    _zz_selectReadFifo_6_40;
  wire       [0:0]    _zz_selectReadFifo_6_41;
  wire       [5:0]    _zz_selectReadFifo_6_42;
  wire       [5:0]    _zz_selectReadFifo_6_43;
  wire       [5:0]    _zz_selectReadFifo_6_44;
  wire       [0:0]    _zz_selectReadFifo_6_45;
  wire       [5:0]    _zz_when_ArraySlice_l165_352;
  wire       [5:0]    _zz_when_ArraySlice_l165_352_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_352_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_352;
  wire       [6:0]    _zz_when_ArraySlice_l166_352_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_352_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_352_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_352_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_352_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_352;
  wire       [6:0]    _zz_when_ArraySlice_l113_352;
  wire       [6:0]    _zz_when_ArraySlice_l113_352_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_352_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_352_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_352_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_352;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_352_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_352_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_352_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_352;
  wire       [6:0]    _zz_when_ArraySlice_l118_352_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_352_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_352_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_352_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_352_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_352_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_352_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_352_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_352_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_353;
  wire       [5:0]    _zz_when_ArraySlice_l165_353_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_353_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_353;
  wire       [5:0]    _zz_when_ArraySlice_l166_353_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_353_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_353_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_353_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_353;
  wire       [6:0]    _zz_when_ArraySlice_l113_353;
  wire       [6:0]    _zz_when_ArraySlice_l113_353_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_353_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_353_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_353_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_353;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_353_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_353_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_353_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_353;
  wire       [6:0]    _zz_when_ArraySlice_l118_353_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_353_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_353_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_353_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_353_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_353_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_353_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_353_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_353_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_353_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_354;
  wire       [5:0]    _zz_when_ArraySlice_l165_354_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_354_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_354;
  wire       [5:0]    _zz_when_ArraySlice_l166_354_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_354_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_354_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_354_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_354;
  wire       [6:0]    _zz_when_ArraySlice_l113_354;
  wire       [6:0]    _zz_when_ArraySlice_l113_354_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_354_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_354_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_354_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_354;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_354_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_354_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_354_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_354;
  wire       [6:0]    _zz_when_ArraySlice_l118_354_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_354_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_354_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_354_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_354_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_354_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_354_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_354_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_354_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_354_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_355;
  wire       [5:0]    _zz_when_ArraySlice_l165_355_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_355_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_355;
  wire       [5:0]    _zz_when_ArraySlice_l166_355_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_355_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_355_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_355_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_355;
  wire       [6:0]    _zz_when_ArraySlice_l113_355;
  wire       [6:0]    _zz_when_ArraySlice_l113_355_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_355_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_355_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_355_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_355;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_355_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_355_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_355_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_355;
  wire       [6:0]    _zz_when_ArraySlice_l118_355_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_355_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_355_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_355_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_355_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_355_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_355_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_355_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_355_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_355_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_356;
  wire       [5:0]    _zz_when_ArraySlice_l165_356_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_356;
  wire       [5:0]    _zz_when_ArraySlice_l166_356_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_356_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_356_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_356;
  wire       [6:0]    _zz_when_ArraySlice_l113_356;
  wire       [6:0]    _zz_when_ArraySlice_l113_356_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_356_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_356_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_356_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_356;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_356_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_356_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_356_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_356;
  wire       [6:0]    _zz_when_ArraySlice_l118_356_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_356_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_356_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_356_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_356_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_356_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_356_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_356_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_356_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_357;
  wire       [5:0]    _zz_when_ArraySlice_l165_357_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_357;
  wire       [4:0]    _zz_when_ArraySlice_l166_357_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_357_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_357_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_357_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_357;
  wire       [6:0]    _zz_when_ArraySlice_l113_357;
  wire       [6:0]    _zz_when_ArraySlice_l113_357_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_357_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_357_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_357_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_357;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_357_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_357_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_357_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_357;
  wire       [6:0]    _zz_when_ArraySlice_l118_357_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_357_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_357_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_357_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_357_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_357_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_357_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_357_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_357_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_358;
  wire       [5:0]    _zz_when_ArraySlice_l165_358_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_358;
  wire       [4:0]    _zz_when_ArraySlice_l166_358_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_358_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_358_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_358_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_358;
  wire       [6:0]    _zz_when_ArraySlice_l113_358;
  wire       [6:0]    _zz_when_ArraySlice_l113_358_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_358_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_358_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_358_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_358;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_358_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_358_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_358_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_358;
  wire       [6:0]    _zz_when_ArraySlice_l118_358_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_358_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_358_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_358_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_358_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_358_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_358_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_358_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_358_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_359;
  wire       [5:0]    _zz_when_ArraySlice_l165_359_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_359;
  wire       [3:0]    _zz_when_ArraySlice_l166_359_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_359_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_359_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_359_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_359;
  wire       [6:0]    _zz_when_ArraySlice_l113_359;
  wire       [6:0]    _zz_when_ArraySlice_l113_359_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_359_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_359_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_359_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_359;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_359_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_359_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_359_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_359;
  wire       [6:0]    _zz_when_ArraySlice_l118_359_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_359_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_359_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_359_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_359_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_359_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_359_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_359_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_359_8;
  wire                _zz_when_ArraySlice_l265_6;
  wire                _zz_when_ArraySlice_l265_6_1;
  wire                _zz_when_ArraySlice_l265_6_2;
  wire                _zz_when_ArraySlice_l265_6_3;
  wire                _zz_when_ArraySlice_l265_6_4;
  wire                _zz_when_ArraySlice_l265_6_5;
  wire       [5:0]    _zz_when_ArraySlice_l268_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l268_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l268_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l268_6_4;
  wire       [5:0]    _zz_when_ArraySlice_l268_6_5;
  wire       [0:0]    _zz_when_ArraySlice_l268_6_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_6_7;
  wire       [5:0]    _zz_selectReadFifo_6_46;
  wire       [0:0]    _zz_selectReadFifo_6_47;
  wire       [12:0]   _zz_when_ArraySlice_l272_6;
  wire       [12:0]   _zz_when_ArraySlice_l272_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l272_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l272_6_3;
  reg        [6:0]    _zz_when_ArraySlice_l276_6;
  wire       [5:0]    _zz_when_ArraySlice_l276_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l276_6_2;
  wire       [12:0]   _zz_when_ArraySlice_l277_6;
  wire       [5:0]    _zz_when_ArraySlice_l277_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l277_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l277_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l277_6_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_43;
  wire       [6:0]    _zz_when_ArraySlice_l95_43;
  wire       [6:0]    _zz_when_ArraySlice_l95_43_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_43_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_43_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_43_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_6;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_6_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_6_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_43;
  wire       [6:0]    _zz_when_ArraySlice_l99_43_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l279_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l279_6_4;
  wire       [5:0]    _zz_selectReadFifo_6_48;
  wire       [5:0]    _zz_selectReadFifo_6_49;
  wire       [5:0]    _zz_selectReadFifo_6_50;
  wire       [0:0]    _zz_selectReadFifo_6_51;
  wire       [5:0]    _zz_selectReadFifo_6_52;
  wire       [5:0]    _zz_selectReadFifo_6_53;
  wire       [5:0]    _zz_selectReadFifo_6_54;
  wire       [0:0]    _zz_selectReadFifo_6_55;
  wire       [5:0]    _zz_when_ArraySlice_l165_360;
  wire       [5:0]    _zz_when_ArraySlice_l165_360_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_360_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_360;
  wire       [6:0]    _zz_when_ArraySlice_l166_360_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_360_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_360_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_360_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_360_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_360;
  wire       [6:0]    _zz_when_ArraySlice_l113_360;
  wire       [6:0]    _zz_when_ArraySlice_l113_360_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_360_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_360_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_360_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_360;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_360_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_360_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_360_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_360;
  wire       [6:0]    _zz_when_ArraySlice_l118_360_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_360_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_360_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_360_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_360_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_360_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_360_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_360_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_360_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_361;
  wire       [5:0]    _zz_when_ArraySlice_l165_361_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_361_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_361;
  wire       [5:0]    _zz_when_ArraySlice_l166_361_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_361_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_361_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_361_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_361;
  wire       [6:0]    _zz_when_ArraySlice_l113_361;
  wire       [6:0]    _zz_when_ArraySlice_l113_361_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_361_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_361_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_361_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_361;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_361_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_361_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_361_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_361;
  wire       [6:0]    _zz_when_ArraySlice_l118_361_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_361_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_361_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_361_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_361_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_361_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_361_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_361_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_361_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_361_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_362;
  wire       [5:0]    _zz_when_ArraySlice_l165_362_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_362_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_362;
  wire       [5:0]    _zz_when_ArraySlice_l166_362_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_362_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_362_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_362_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_362;
  wire       [6:0]    _zz_when_ArraySlice_l113_362;
  wire       [6:0]    _zz_when_ArraySlice_l113_362_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_362_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_362_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_362_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_362;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_362_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_362_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_362_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_362;
  wire       [6:0]    _zz_when_ArraySlice_l118_362_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_362_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_362_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_362_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_362_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_362_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_362_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_362_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_362_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_362_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_363;
  wire       [5:0]    _zz_when_ArraySlice_l165_363_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_363_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_363;
  wire       [5:0]    _zz_when_ArraySlice_l166_363_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_363_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_363_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_363_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_363;
  wire       [6:0]    _zz_when_ArraySlice_l113_363;
  wire       [6:0]    _zz_when_ArraySlice_l113_363_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_363_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_363_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_363_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_363;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_363_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_363_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_363_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_363;
  wire       [6:0]    _zz_when_ArraySlice_l118_363_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_363_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_363_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_363_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_363_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_363_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_363_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_363_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_363_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_363_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_364;
  wire       [5:0]    _zz_when_ArraySlice_l165_364_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_364;
  wire       [5:0]    _zz_when_ArraySlice_l166_364_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_364_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_364_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_364;
  wire       [6:0]    _zz_when_ArraySlice_l113_364;
  wire       [6:0]    _zz_when_ArraySlice_l113_364_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_364_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_364_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_364_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_364;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_364_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_364_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_364_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_364;
  wire       [6:0]    _zz_when_ArraySlice_l118_364_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_364_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_364_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_364_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_364_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_364_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_364_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_364_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_364_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_365;
  wire       [5:0]    _zz_when_ArraySlice_l165_365_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_365;
  wire       [4:0]    _zz_when_ArraySlice_l166_365_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_365_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_365_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_365_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_365;
  wire       [6:0]    _zz_when_ArraySlice_l113_365;
  wire       [6:0]    _zz_when_ArraySlice_l113_365_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_365_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_365_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_365_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_365;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_365_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_365_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_365_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_365;
  wire       [6:0]    _zz_when_ArraySlice_l118_365_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_365_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_365_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_365_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_365_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_365_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_365_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_365_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_365_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_366;
  wire       [5:0]    _zz_when_ArraySlice_l165_366_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_366;
  wire       [4:0]    _zz_when_ArraySlice_l166_366_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_366_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_366_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_366_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_366;
  wire       [6:0]    _zz_when_ArraySlice_l113_366;
  wire       [6:0]    _zz_when_ArraySlice_l113_366_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_366_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_366_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_366_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_366;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_366_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_366_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_366_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_366;
  wire       [6:0]    _zz_when_ArraySlice_l118_366_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_366_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_366_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_366_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_366_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_366_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_366_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_366_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_366_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_367;
  wire       [5:0]    _zz_when_ArraySlice_l165_367_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_367;
  wire       [3:0]    _zz_when_ArraySlice_l166_367_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_367_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_367_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_367_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_367;
  wire       [6:0]    _zz_when_ArraySlice_l113_367;
  wire       [6:0]    _zz_when_ArraySlice_l113_367_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_367_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_367_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_367_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_367;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_367_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_367_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_367_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_367;
  wire       [6:0]    _zz_when_ArraySlice_l118_367_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_367_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_367_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_367_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_367_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_367_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_367_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_367_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_367_8;
  wire                _zz_when_ArraySlice_l285_6;
  wire                _zz_when_ArraySlice_l285_6_1;
  wire                _zz_when_ArraySlice_l285_6_2;
  wire                _zz_when_ArraySlice_l285_6_3;
  wire                _zz_when_ArraySlice_l285_6_4;
  wire                _zz_when_ArraySlice_l285_6_5;
  wire       [5:0]    _zz_when_ArraySlice_l288_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l288_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l288_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l288_6_4;
  wire       [5:0]    _zz_when_ArraySlice_l288_6_5;
  wire       [0:0]    _zz_when_ArraySlice_l288_6_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_6_7;
  wire       [5:0]    _zz_selectReadFifo_6_56;
  wire       [0:0]    _zz_selectReadFifo_6_57;
  wire       [12:0]   _zz_when_ArraySlice_l292_6;
  wire       [12:0]   _zz_when_ArraySlice_l292_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l292_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l292_6_3;
  wire       [12:0]   _zz_when_ArraySlice_l303_6;
  wire       [5:0]    _zz_when_ArraySlice_l303_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l303_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l303_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l303_6_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_44;
  wire       [6:0]    _zz_when_ArraySlice_l95_44;
  wire       [6:0]    _zz_when_ArraySlice_l95_44_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_44_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_44_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_44_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_6;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_6_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_6_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_44;
  wire       [6:0]    _zz_when_ArraySlice_l99_44_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l304_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l304_6_4;
  wire       [5:0]    _zz_selectReadFifo_6_58;
  wire       [5:0]    _zz_selectReadFifo_6_59;
  wire       [5:0]    _zz_selectReadFifo_6_60;
  wire       [0:0]    _zz_selectReadFifo_6_61;
  wire       [5:0]    _zz_when_ArraySlice_l165_368;
  wire       [5:0]    _zz_when_ArraySlice_l165_368_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_368_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_368;
  wire       [6:0]    _zz_when_ArraySlice_l166_368_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_368_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_368_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_368_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_368_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_368;
  wire       [6:0]    _zz_when_ArraySlice_l113_368;
  wire       [6:0]    _zz_when_ArraySlice_l113_368_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_368_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_368_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_368_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_368;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_368_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_368_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_368_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_368;
  wire       [6:0]    _zz_when_ArraySlice_l118_368_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_368_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_368_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_368_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_368_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_368_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_368_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_368_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_368_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_369;
  wire       [5:0]    _zz_when_ArraySlice_l165_369_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_369_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_369;
  wire       [5:0]    _zz_when_ArraySlice_l166_369_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_369_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_369_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_369_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_369;
  wire       [6:0]    _zz_when_ArraySlice_l113_369;
  wire       [6:0]    _zz_when_ArraySlice_l113_369_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_369_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_369_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_369_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_369;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_369_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_369_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_369_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_369;
  wire       [6:0]    _zz_when_ArraySlice_l118_369_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_369_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_369_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_369_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_369_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_369_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_369_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_369_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_369_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_369_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_370;
  wire       [5:0]    _zz_when_ArraySlice_l165_370_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_370_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_370;
  wire       [5:0]    _zz_when_ArraySlice_l166_370_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_370_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_370_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_370_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_370;
  wire       [6:0]    _zz_when_ArraySlice_l113_370;
  wire       [6:0]    _zz_when_ArraySlice_l113_370_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_370_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_370_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_370_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_370;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_370_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_370_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_370_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_370;
  wire       [6:0]    _zz_when_ArraySlice_l118_370_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_370_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_370_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_370_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_370_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_370_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_370_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_370_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_370_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_370_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_371;
  wire       [5:0]    _zz_when_ArraySlice_l165_371_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_371_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_371;
  wire       [5:0]    _zz_when_ArraySlice_l166_371_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_371_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_371_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_371_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_371;
  wire       [6:0]    _zz_when_ArraySlice_l113_371;
  wire       [6:0]    _zz_when_ArraySlice_l113_371_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_371_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_371_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_371_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_371;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_371_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_371_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_371_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_371;
  wire       [6:0]    _zz_when_ArraySlice_l118_371_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_371_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_371_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_371_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_371_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_371_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_371_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_371_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_371_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_371_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_372;
  wire       [5:0]    _zz_when_ArraySlice_l165_372_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_372;
  wire       [5:0]    _zz_when_ArraySlice_l166_372_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_372_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_372_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_372;
  wire       [6:0]    _zz_when_ArraySlice_l113_372;
  wire       [6:0]    _zz_when_ArraySlice_l113_372_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_372_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_372_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_372_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_372;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_372_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_372_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_372_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_372;
  wire       [6:0]    _zz_when_ArraySlice_l118_372_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_372_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_372_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_372_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_372_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_372_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_372_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_372_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_372_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_373;
  wire       [5:0]    _zz_when_ArraySlice_l165_373_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_373;
  wire       [4:0]    _zz_when_ArraySlice_l166_373_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_373_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_373_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_373_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_373;
  wire       [6:0]    _zz_when_ArraySlice_l113_373;
  wire       [6:0]    _zz_when_ArraySlice_l113_373_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_373_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_373_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_373_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_373;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_373_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_373_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_373_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_373;
  wire       [6:0]    _zz_when_ArraySlice_l118_373_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_373_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_373_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_373_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_373_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_373_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_373_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_373_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_373_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_374;
  wire       [5:0]    _zz_when_ArraySlice_l165_374_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_374;
  wire       [4:0]    _zz_when_ArraySlice_l166_374_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_374_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_374_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_374_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_374;
  wire       [6:0]    _zz_when_ArraySlice_l113_374;
  wire       [6:0]    _zz_when_ArraySlice_l113_374_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_374_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_374_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_374_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_374;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_374_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_374_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_374_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_374;
  wire       [6:0]    _zz_when_ArraySlice_l118_374_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_374_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_374_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_374_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_374_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_374_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_374_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_374_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_374_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_375;
  wire       [5:0]    _zz_when_ArraySlice_l165_375_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_375;
  wire       [3:0]    _zz_when_ArraySlice_l166_375_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_375_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_375_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_375_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_375;
  wire       [6:0]    _zz_when_ArraySlice_l113_375;
  wire       [6:0]    _zz_when_ArraySlice_l113_375_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_375_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_375_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_375_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_375;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_375_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_375_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_375_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_375;
  wire       [6:0]    _zz_when_ArraySlice_l118_375_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_375_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_375_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_375_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_375_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_375_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_375_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_375_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_375_8;
  wire                _zz_when_ArraySlice_l311_6;
  wire                _zz_when_ArraySlice_l311_6_1;
  wire                _zz_when_ArraySlice_l311_6_2;
  wire                _zz_when_ArraySlice_l311_6_3;
  wire                _zz_when_ArraySlice_l311_6_4;
  wire                _zz_when_ArraySlice_l311_6_5;
  wire       [5:0]    _zz_selectReadFifo_6_62;
  wire       [0:0]    _zz_selectReadFifo_6_63;
  wire       [12:0]   _zz_when_ArraySlice_l315_6;
  wire       [12:0]   _zz_when_ArraySlice_l315_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l315_6_2;
  wire       [0:0]    _zz_when_ArraySlice_l315_6_3;
  wire       [5:0]    _zz_when_ArraySlice_l301_6;
  wire       [5:0]    _zz_when_ArraySlice_l301_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l322_6;
  wire       [5:0]    _zz_when_ArraySlice_l322_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l322_6_2;
  wire       [5:0]    _zz_when_ArraySlice_l322_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l322_6_4;
  wire       [5:0]    _zz_when_ArraySlice_l240_7;
  wire       [5:0]    _zz_when_ArraySlice_l240_7_1;
  reg        [6:0]    _zz_when_ArraySlice_l241_7;
  wire       [5:0]    _zz_when_ArraySlice_l241_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l241_7_2;
  wire       [5:0]    _zz__zz_outputStreamArrayData_7_valid_1;
  reg                 _zz_outputStreamArrayData_7_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_7_payload_1;
  wire       [6:0]    _zz_when_ArraySlice_l247_7;
  wire       [0:0]    _zz_when_ArraySlice_l247_7_1;
  reg        [6:0]    _zz_when_ArraySlice_l247_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l247_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l247_7_4;
  wire       [12:0]   _zz_when_ArraySlice_l248_7;
  wire       [5:0]    _zz_when_ArraySlice_l248_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l248_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l248_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l248_7_4;
  wire       [5:0]    _zz_selectReadFifo_7_32;
  wire       [5:0]    _zz_selectReadFifo_7_33;
  wire       [5:0]    _zz_selectReadFifo_7_34;
  wire       [0:0]    _zz_selectReadFifo_7_35;
  wire       [5:0]    _zz_selectReadFifo_7_36;
  wire       [0:0]    _zz_selectReadFifo_7_37;
  wire       [12:0]   _zz_when_ArraySlice_l251_7;
  wire       [12:0]   _zz_when_ArraySlice_l251_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l251_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l251_7_3;
  reg        [6:0]    _zz_when_ArraySlice_l256_7;
  wire       [5:0]    _zz_when_ArraySlice_l256_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l256_7_2;
  wire       [6:0]    _zz_when_ArraySlice_l256_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l256_7_4;
  wire       [12:0]   _zz_when_ArraySlice_l257_7;
  wire       [5:0]    _zz_when_ArraySlice_l257_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l257_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l257_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l257_7_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_45;
  wire       [6:0]    _zz_when_ArraySlice_l95_45;
  wire       [6:0]    _zz_when_ArraySlice_l95_45_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_45_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_45_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_45_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_7;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_7_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_7_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l259_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_45;
  wire       [6:0]    _zz_when_ArraySlice_l99_45_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l259_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l259_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l259_7_4;
  wire       [5:0]    _zz_selectReadFifo_7_38;
  wire       [5:0]    _zz_selectReadFifo_7_39;
  wire       [5:0]    _zz_selectReadFifo_7_40;
  wire       [0:0]    _zz_selectReadFifo_7_41;
  wire       [5:0]    _zz_selectReadFifo_7_42;
  wire       [5:0]    _zz_selectReadFifo_7_43;
  wire       [5:0]    _zz_selectReadFifo_7_44;
  wire       [0:0]    _zz_selectReadFifo_7_45;
  wire       [5:0]    _zz_when_ArraySlice_l165_376;
  wire       [5:0]    _zz_when_ArraySlice_l165_376_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_376_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_376;
  wire       [6:0]    _zz_when_ArraySlice_l166_376_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_376_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_376_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_376_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_376_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_376;
  wire       [6:0]    _zz_when_ArraySlice_l113_376;
  wire       [6:0]    _zz_when_ArraySlice_l113_376_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_376_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_376_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_376_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_376;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_376_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_376_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_376_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_376;
  wire       [6:0]    _zz_when_ArraySlice_l118_376_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_376_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_376_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_376_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_376_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_376_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_376_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_376_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_376_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_377;
  wire       [5:0]    _zz_when_ArraySlice_l165_377_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_377_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_377;
  wire       [5:0]    _zz_when_ArraySlice_l166_377_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_377_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_377_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_377_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_377;
  wire       [6:0]    _zz_when_ArraySlice_l113_377;
  wire       [6:0]    _zz_when_ArraySlice_l113_377_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_377_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_377_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_377_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_377;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_377_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_377_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_377_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_377;
  wire       [6:0]    _zz_when_ArraySlice_l118_377_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_377_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_377_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_377_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_377_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_377_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_377_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_377_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_377_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_377_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_378;
  wire       [5:0]    _zz_when_ArraySlice_l165_378_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_378_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_378;
  wire       [5:0]    _zz_when_ArraySlice_l166_378_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_378_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_378_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_378_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_378;
  wire       [6:0]    _zz_when_ArraySlice_l113_378;
  wire       [6:0]    _zz_when_ArraySlice_l113_378_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_378_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_378_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_378_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_378;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_378_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_378_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_378_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_378;
  wire       [6:0]    _zz_when_ArraySlice_l118_378_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_378_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_378_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_378_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_378_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_378_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_378_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_378_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_378_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_378_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_379;
  wire       [5:0]    _zz_when_ArraySlice_l165_379_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_379_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_379;
  wire       [5:0]    _zz_when_ArraySlice_l166_379_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_379_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_379_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_379_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_379;
  wire       [6:0]    _zz_when_ArraySlice_l113_379;
  wire       [6:0]    _zz_when_ArraySlice_l113_379_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_379_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_379_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_379_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_379;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_379_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_379_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_379_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_379;
  wire       [6:0]    _zz_when_ArraySlice_l118_379_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_379_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_379_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_379_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_379_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_379_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_379_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_379_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_379_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_379_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_380;
  wire       [5:0]    _zz_when_ArraySlice_l165_380_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_380;
  wire       [5:0]    _zz_when_ArraySlice_l166_380_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_380_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_380_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_380;
  wire       [6:0]    _zz_when_ArraySlice_l113_380;
  wire       [6:0]    _zz_when_ArraySlice_l113_380_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_380_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_380_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_380_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_380;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_380_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_380_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_380_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_380;
  wire       [6:0]    _zz_when_ArraySlice_l118_380_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_380_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_380_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_380_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_380_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_380_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_380_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_380_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_380_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_381;
  wire       [5:0]    _zz_when_ArraySlice_l165_381_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_381;
  wire       [4:0]    _zz_when_ArraySlice_l166_381_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_381_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_381_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_381_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_381;
  wire       [6:0]    _zz_when_ArraySlice_l113_381;
  wire       [6:0]    _zz_when_ArraySlice_l113_381_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_381_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_381_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_381_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_381;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_381_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_381_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_381_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_381;
  wire       [6:0]    _zz_when_ArraySlice_l118_381_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_381_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_381_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_381_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_381_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_381_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_381_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_381_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_381_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_382;
  wire       [5:0]    _zz_when_ArraySlice_l165_382_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_382;
  wire       [4:0]    _zz_when_ArraySlice_l166_382_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_382_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_382_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_382_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_382;
  wire       [6:0]    _zz_when_ArraySlice_l113_382;
  wire       [6:0]    _zz_when_ArraySlice_l113_382_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_382_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_382_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_382_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_382;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_382_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_382_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_382_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_382;
  wire       [6:0]    _zz_when_ArraySlice_l118_382_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_382_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_382_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_382_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_382_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_382_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_382_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_382_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_382_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_383;
  wire       [5:0]    _zz_when_ArraySlice_l165_383_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_383;
  wire       [3:0]    _zz_when_ArraySlice_l166_383_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_383_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_383_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_383_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_383;
  wire       [6:0]    _zz_when_ArraySlice_l113_383;
  wire       [6:0]    _zz_when_ArraySlice_l113_383_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_383_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_383_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_383_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_383;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_383_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_383_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_383_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_383;
  wire       [6:0]    _zz_when_ArraySlice_l118_383_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_383_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_383_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_383_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_383_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_383_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_383_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_383_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_383_8;
  wire                _zz_when_ArraySlice_l265_7;
  wire                _zz_when_ArraySlice_l265_7_1;
  wire                _zz_when_ArraySlice_l265_7_2;
  wire                _zz_when_ArraySlice_l265_7_3;
  wire                _zz_when_ArraySlice_l265_7_4;
  wire                _zz_when_ArraySlice_l265_7_5;
  wire       [5:0]    _zz_when_ArraySlice_l268_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l268_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l268_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l268_7_4;
  wire       [5:0]    _zz_when_ArraySlice_l268_7_5;
  wire       [0:0]    _zz_when_ArraySlice_l268_7_6;
  wire       [5:0]    _zz_when_ArraySlice_l268_7_7;
  wire       [5:0]    _zz_selectReadFifo_7_46;
  wire       [0:0]    _zz_selectReadFifo_7_47;
  wire       [12:0]   _zz_when_ArraySlice_l272_7;
  wire       [12:0]   _zz_when_ArraySlice_l272_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l272_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l272_7_3;
  reg        [6:0]    _zz_when_ArraySlice_l276_7;
  wire       [5:0]    _zz_when_ArraySlice_l276_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l276_7_2;
  wire       [12:0]   _zz_when_ArraySlice_l277_7;
  wire       [5:0]    _zz_when_ArraySlice_l277_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l277_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l277_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l277_7_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_46;
  wire       [6:0]    _zz_when_ArraySlice_l95_46;
  wire       [6:0]    _zz_when_ArraySlice_l95_46_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_46_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_46_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_46_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_7;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_7_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_7_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l279_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_46;
  wire       [6:0]    _zz_when_ArraySlice_l99_46_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l279_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l279_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l279_7_4;
  wire       [5:0]    _zz_selectReadFifo_7_48;
  wire       [5:0]    _zz_selectReadFifo_7_49;
  wire       [5:0]    _zz_selectReadFifo_7_50;
  wire       [0:0]    _zz_selectReadFifo_7_51;
  wire       [5:0]    _zz_selectReadFifo_7_52;
  wire       [5:0]    _zz_selectReadFifo_7_53;
  wire       [5:0]    _zz_selectReadFifo_7_54;
  wire       [0:0]    _zz_selectReadFifo_7_55;
  wire       [5:0]    _zz_when_ArraySlice_l165_384;
  wire       [5:0]    _zz_when_ArraySlice_l165_384_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_384_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_384;
  wire       [6:0]    _zz_when_ArraySlice_l166_384_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_384_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_384_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_384_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_384_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_384;
  wire       [6:0]    _zz_when_ArraySlice_l113_384;
  wire       [6:0]    _zz_when_ArraySlice_l113_384_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_384_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_384_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_384_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_384;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_384_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_384_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_384_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_384;
  wire       [6:0]    _zz_when_ArraySlice_l118_384_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_384_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_384_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_384_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_384_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_384_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_384_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_384_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_384_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_385;
  wire       [5:0]    _zz_when_ArraySlice_l165_385_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_385_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_385;
  wire       [5:0]    _zz_when_ArraySlice_l166_385_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_385_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_385_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_385_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_385;
  wire       [6:0]    _zz_when_ArraySlice_l113_385;
  wire       [6:0]    _zz_when_ArraySlice_l113_385_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_385_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_385_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_385_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_385;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_385_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_385_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_385_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_385;
  wire       [6:0]    _zz_when_ArraySlice_l118_385_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_385_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_385_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_385_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_385_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_385_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_385_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_385_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_385_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_385_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_386;
  wire       [5:0]    _zz_when_ArraySlice_l165_386_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_386_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_386;
  wire       [5:0]    _zz_when_ArraySlice_l166_386_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_386_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_386_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_386_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_386;
  wire       [6:0]    _zz_when_ArraySlice_l113_386;
  wire       [6:0]    _zz_when_ArraySlice_l113_386_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_386_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_386_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_386_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_386;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_386_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_386_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_386_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_386;
  wire       [6:0]    _zz_when_ArraySlice_l118_386_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_386_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_386_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_386_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_386_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_386_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_386_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_386_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_386_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_386_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_387;
  wire       [5:0]    _zz_when_ArraySlice_l165_387_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_387_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_387;
  wire       [5:0]    _zz_when_ArraySlice_l166_387_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_387_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_387_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_387_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_387;
  wire       [6:0]    _zz_when_ArraySlice_l113_387;
  wire       [6:0]    _zz_when_ArraySlice_l113_387_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_387_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_387_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_387_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_387;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_387_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_387_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_387_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_387;
  wire       [6:0]    _zz_when_ArraySlice_l118_387_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_387_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_387_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_387_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_387_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_387_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_387_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_387_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_387_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_387_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_388;
  wire       [5:0]    _zz_when_ArraySlice_l165_388_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_388;
  wire       [5:0]    _zz_when_ArraySlice_l166_388_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_388_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_388_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_388;
  wire       [6:0]    _zz_when_ArraySlice_l113_388;
  wire       [6:0]    _zz_when_ArraySlice_l113_388_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_388_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_388_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_388_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_388;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_388_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_388_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_388_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_388;
  wire       [6:0]    _zz_when_ArraySlice_l118_388_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_388_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_388_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_388_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_388_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_388_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_388_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_388_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_388_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_389;
  wire       [5:0]    _zz_when_ArraySlice_l165_389_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_389;
  wire       [4:0]    _zz_when_ArraySlice_l166_389_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_389_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_389_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_389_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_389;
  wire       [6:0]    _zz_when_ArraySlice_l113_389;
  wire       [6:0]    _zz_when_ArraySlice_l113_389_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_389_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_389_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_389_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_389;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_389_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_389_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_389_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_389;
  wire       [6:0]    _zz_when_ArraySlice_l118_389_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_389_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_389_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_389_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_389_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_389_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_389_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_389_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_389_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_390;
  wire       [5:0]    _zz_when_ArraySlice_l165_390_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_390;
  wire       [4:0]    _zz_when_ArraySlice_l166_390_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_390_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_390_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_390_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_390;
  wire       [6:0]    _zz_when_ArraySlice_l113_390;
  wire       [6:0]    _zz_when_ArraySlice_l113_390_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_390_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_390_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_390_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_390;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_390_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_390_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_390_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_390;
  wire       [6:0]    _zz_when_ArraySlice_l118_390_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_390_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_390_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_390_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_390_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_390_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_390_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_390_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_390_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_391;
  wire       [5:0]    _zz_when_ArraySlice_l165_391_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_391;
  wire       [3:0]    _zz_when_ArraySlice_l166_391_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_391_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_391_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_391_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_391;
  wire       [6:0]    _zz_when_ArraySlice_l113_391;
  wire       [6:0]    _zz_when_ArraySlice_l113_391_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_391_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_391_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_391_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_391;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_391_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_391_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_391_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_391;
  wire       [6:0]    _zz_when_ArraySlice_l118_391_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_391_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_391_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_391_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_391_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_391_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_391_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_391_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_391_8;
  wire                _zz_when_ArraySlice_l285_7;
  wire                _zz_when_ArraySlice_l285_7_1;
  wire                _zz_when_ArraySlice_l285_7_2;
  wire                _zz_when_ArraySlice_l285_7_3;
  wire                _zz_when_ArraySlice_l285_7_4;
  wire                _zz_when_ArraySlice_l285_7_5;
  wire       [5:0]    _zz_when_ArraySlice_l288_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l288_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l288_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l288_7_4;
  wire       [5:0]    _zz_when_ArraySlice_l288_7_5;
  wire       [0:0]    _zz_when_ArraySlice_l288_7_6;
  wire       [5:0]    _zz_when_ArraySlice_l288_7_7;
  wire       [5:0]    _zz_selectReadFifo_7_56;
  wire       [0:0]    _zz_selectReadFifo_7_57;
  wire       [12:0]   _zz_when_ArraySlice_l292_7;
  wire       [12:0]   _zz_when_ArraySlice_l292_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l292_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l292_7_3;
  wire       [12:0]   _zz_when_ArraySlice_l303_7;
  wire       [5:0]    _zz_when_ArraySlice_l303_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l303_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l303_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l303_7_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l94_47;
  wire       [6:0]    _zz_when_ArraySlice_l95_47;
  wire       [6:0]    _zz_when_ArraySlice_l95_47_1;
  wire       [6:0]    _zz_when_ArraySlice_l95_47_2;
  wire       [6:0]    _zz_when_ArraySlice_l95_47_3;
  wire       [6:0]    _zz_when_ArraySlice_l95_47_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_7;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_7_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_7_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l304_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l99_47;
  wire       [6:0]    _zz_when_ArraySlice_l99_47_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l304_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l304_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l304_7_4;
  wire       [5:0]    _zz_selectReadFifo_7_58;
  wire       [5:0]    _zz_selectReadFifo_7_59;
  wire       [5:0]    _zz_selectReadFifo_7_60;
  wire       [0:0]    _zz_selectReadFifo_7_61;
  wire       [5:0]    _zz_when_ArraySlice_l165_392;
  wire       [5:0]    _zz_when_ArraySlice_l165_392_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_392_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_392;
  wire       [6:0]    _zz_when_ArraySlice_l166_392_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_392_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_392_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_392_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_392_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_392;
  wire       [6:0]    _zz_when_ArraySlice_l113_392;
  wire       [6:0]    _zz_when_ArraySlice_l113_392_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_392_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_392_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_392_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_392;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_392_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_392_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_392_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_392;
  wire       [6:0]    _zz_when_ArraySlice_l118_392_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_392_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_392_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_392_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_392_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_392_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_392_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_392_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_392_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_393;
  wire       [5:0]    _zz_when_ArraySlice_l165_393_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_393_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_393;
  wire       [5:0]    _zz_when_ArraySlice_l166_393_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_393_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_393_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_393_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_393;
  wire       [6:0]    _zz_when_ArraySlice_l113_393;
  wire       [6:0]    _zz_when_ArraySlice_l113_393_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_393_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_393_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_393_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_393;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_393_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_393_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_393_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_393;
  wire       [6:0]    _zz_when_ArraySlice_l118_393_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_393_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_393_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_393_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_393_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_393_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_393_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_393_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_393_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_393_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_394;
  wire       [5:0]    _zz_when_ArraySlice_l165_394_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_394_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_394;
  wire       [5:0]    _zz_when_ArraySlice_l166_394_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_394_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_394_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_394_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_394;
  wire       [6:0]    _zz_when_ArraySlice_l113_394;
  wire       [6:0]    _zz_when_ArraySlice_l113_394_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_394_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_394_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_394_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_394;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_394_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_394_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_394_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_394;
  wire       [6:0]    _zz_when_ArraySlice_l118_394_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_394_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_394_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_394_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_394_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_394_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_394_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_394_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_394_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_394_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_395;
  wire       [5:0]    _zz_when_ArraySlice_l165_395_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_395_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_395;
  wire       [5:0]    _zz_when_ArraySlice_l166_395_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_395_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_395_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_395_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_395;
  wire       [6:0]    _zz_when_ArraySlice_l113_395;
  wire       [6:0]    _zz_when_ArraySlice_l113_395_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_395_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_395_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_395_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_395;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_395_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_395_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_395_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_395;
  wire       [6:0]    _zz_when_ArraySlice_l118_395_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_395_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_395_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_395_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_395_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_395_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_395_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_395_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_395_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_395_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_396;
  wire       [5:0]    _zz_when_ArraySlice_l165_396_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_396;
  wire       [5:0]    _zz_when_ArraySlice_l166_396_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_396_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_396_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_396;
  wire       [6:0]    _zz_when_ArraySlice_l113_396;
  wire       [6:0]    _zz_when_ArraySlice_l113_396_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_396_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_396_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_396_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_396;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_396_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_396_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_396_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_396;
  wire       [6:0]    _zz_when_ArraySlice_l118_396_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_396_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_396_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_396_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_396_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_396_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_396_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_396_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_396_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_397;
  wire       [5:0]    _zz_when_ArraySlice_l165_397_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_397;
  wire       [4:0]    _zz_when_ArraySlice_l166_397_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_397_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_397_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_397_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_397;
  wire       [6:0]    _zz_when_ArraySlice_l113_397;
  wire       [6:0]    _zz_when_ArraySlice_l113_397_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_397_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_397_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_397_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_397;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_397_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_397_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_397_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_397;
  wire       [6:0]    _zz_when_ArraySlice_l118_397_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_397_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_397_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_397_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_397_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_397_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_397_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_397_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_397_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_398;
  wire       [5:0]    _zz_when_ArraySlice_l165_398_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_398;
  wire       [4:0]    _zz_when_ArraySlice_l166_398_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_398_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_398_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_398_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_398;
  wire       [6:0]    _zz_when_ArraySlice_l113_398;
  wire       [6:0]    _zz_when_ArraySlice_l113_398_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_398_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_398_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_398_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_398;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_398_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_398_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_398_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_398;
  wire       [6:0]    _zz_when_ArraySlice_l118_398_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_398_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_398_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_398_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_398_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_398_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_398_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_398_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_398_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_399;
  wire       [5:0]    _zz_when_ArraySlice_l165_399_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_399;
  wire       [3:0]    _zz_when_ArraySlice_l166_399_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_399_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_399_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_399_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_399;
  wire       [6:0]    _zz_when_ArraySlice_l113_399;
  wire       [6:0]    _zz_when_ArraySlice_l113_399_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_399_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_399_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_399_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_399;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_399_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_399_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_399_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_399;
  wire       [6:0]    _zz_when_ArraySlice_l118_399_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_399_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_399_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_399_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_399_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_399_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_399_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_399_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_399_8;
  wire                _zz_when_ArraySlice_l311_7;
  wire                _zz_when_ArraySlice_l311_7_1;
  wire                _zz_when_ArraySlice_l311_7_2;
  wire                _zz_when_ArraySlice_l311_7_3;
  wire                _zz_when_ArraySlice_l311_7_4;
  wire                _zz_when_ArraySlice_l311_7_5;
  wire       [5:0]    _zz_selectReadFifo_7_62;
  wire       [0:0]    _zz_selectReadFifo_7_63;
  wire       [12:0]   _zz_when_ArraySlice_l315_7;
  wire       [12:0]   _zz_when_ArraySlice_l315_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l315_7_2;
  wire       [0:0]    _zz_when_ArraySlice_l315_7_3;
  wire       [5:0]    _zz_when_ArraySlice_l301_7;
  wire       [5:0]    _zz_when_ArraySlice_l301_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l322_7;
  wire       [5:0]    _zz_when_ArraySlice_l322_7_1;
  wire       [5:0]    _zz_when_ArraySlice_l322_7_2;
  wire       [5:0]    _zz_when_ArraySlice_l322_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l322_7_4;
  wire       [5:0]    _zz_when_ArraySlice_l189;
  wire       [5:0]    _zz_when_ArraySlice_l189_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_1_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_1_2;
  wire       [5:0]    _zz_when_ArraySlice_l189_2;
  wire       [5:0]    _zz_when_ArraySlice_l189_2_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_3;
  wire       [5:0]    _zz_when_ArraySlice_l189_3_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_4;
  wire       [5:0]    _zz_when_ArraySlice_l189_4_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_5;
  wire       [5:0]    _zz_when_ArraySlice_l189_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_6;
  wire       [5:0]    _zz_when_ArraySlice_l189_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_7;
  wire       [5:0]    _zz_when_ArraySlice_l189_7_1;
  wire                _zz_when_ArraySlice_l333_8;
  wire                _zz_when_ArraySlice_l333_9;
  reg        [6:0]    _zz_when_ArraySlice_l334;
  wire       [6:0]    _zz_when_ArraySlice_l334_1;
  reg                 _zz_inputStreamArrayData_ready_1;
  reg        [6:0]    _zz_when_ArraySlice_l338;
  wire       [6:0]    _zz_when_ArraySlice_l338_1;
  wire       [5:0]    _zz_when_ArraySlice_l338_2;
  wire       [5:0]    _zz_when_ArraySlice_l338_3;
  wire       [0:0]    _zz_when_ArraySlice_l338_4;
  wire       [5:0]    _zz_when_ArraySlice_l339;
  wire       [5:0]    _zz_when_ArraySlice_l339_1;
  wire       [0:0]    _zz_when_ArraySlice_l339_2;
  wire       [5:0]    _zz_selectWriteFifo_2;
  wire       [0:0]    _zz_selectWriteFifo_3;
  wire       [5:0]    _zz_when_ArraySlice_l165_400;
  wire       [5:0]    _zz_when_ArraySlice_l165_400_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_400_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_400;
  wire       [6:0]    _zz_when_ArraySlice_l166_400_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_400_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_400_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_400_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_400_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_400;
  wire       [6:0]    _zz_when_ArraySlice_l113_400;
  wire       [6:0]    _zz_when_ArraySlice_l113_400_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_400_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_400_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_400_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_400;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_400_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_400_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_400_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_400;
  wire       [6:0]    _zz_when_ArraySlice_l118_400_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_400_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_400_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_400_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_400_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_400_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_400_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_400_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_400_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_401;
  wire       [5:0]    _zz_when_ArraySlice_l165_401_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_401_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_401;
  wire       [5:0]    _zz_when_ArraySlice_l166_401_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_401_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_401_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_401_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_401;
  wire       [6:0]    _zz_when_ArraySlice_l113_401;
  wire       [6:0]    _zz_when_ArraySlice_l113_401_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_401_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_401_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_401_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_401;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_401_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_401_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_401_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_401;
  wire       [6:0]    _zz_when_ArraySlice_l118_401_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_401_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_401_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_401_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_401_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_401_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_401_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_401_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_401_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_401_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_402;
  wire       [5:0]    _zz_when_ArraySlice_l165_402_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_402_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_402;
  wire       [5:0]    _zz_when_ArraySlice_l166_402_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_402_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_402_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_402_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_402;
  wire       [6:0]    _zz_when_ArraySlice_l113_402;
  wire       [6:0]    _zz_when_ArraySlice_l113_402_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_402_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_402_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_402_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_402;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_402_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_402_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_402_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_402;
  wire       [6:0]    _zz_when_ArraySlice_l118_402_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_402_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_402_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_402_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_402_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_402_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_402_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_402_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_402_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_402_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_403;
  wire       [5:0]    _zz_when_ArraySlice_l165_403_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_403_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_403;
  wire       [5:0]    _zz_when_ArraySlice_l166_403_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_403_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_403_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_403_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_403;
  wire       [6:0]    _zz_when_ArraySlice_l113_403;
  wire       [6:0]    _zz_when_ArraySlice_l113_403_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_403_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_403_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_403_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_403;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_403_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_403_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_403_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_403;
  wire       [6:0]    _zz_when_ArraySlice_l118_403_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_403_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_403_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_403_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_403_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_403_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_403_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_403_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_403_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_403_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_404;
  wire       [5:0]    _zz_when_ArraySlice_l165_404_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_404;
  wire       [5:0]    _zz_when_ArraySlice_l166_404_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_404_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_404_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_404;
  wire       [6:0]    _zz_when_ArraySlice_l113_404;
  wire       [6:0]    _zz_when_ArraySlice_l113_404_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_404_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_404_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_404_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_404;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_404_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_404_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_404_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_404;
  wire       [6:0]    _zz_when_ArraySlice_l118_404_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_404_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_404_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_404_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_404_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_404_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_404_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_404_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_404_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_405;
  wire       [5:0]    _zz_when_ArraySlice_l165_405_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_405;
  wire       [4:0]    _zz_when_ArraySlice_l166_405_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_405_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_405_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_405_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_405;
  wire       [6:0]    _zz_when_ArraySlice_l113_405;
  wire       [6:0]    _zz_when_ArraySlice_l113_405_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_405_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_405_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_405_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_405;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_405_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_405_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_405_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_405;
  wire       [6:0]    _zz_when_ArraySlice_l118_405_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_405_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_405_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_405_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_405_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_405_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_405_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_405_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_405_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_406;
  wire       [5:0]    _zz_when_ArraySlice_l165_406_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_406;
  wire       [4:0]    _zz_when_ArraySlice_l166_406_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_406_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_406_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_406_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_406;
  wire       [6:0]    _zz_when_ArraySlice_l113_406;
  wire       [6:0]    _zz_when_ArraySlice_l113_406_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_406_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_406_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_406_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_406;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_406_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_406_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_406_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_406;
  wire       [6:0]    _zz_when_ArraySlice_l118_406_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_406_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_406_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_406_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_406_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_406_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_406_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_406_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_406_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_407;
  wire       [5:0]    _zz_when_ArraySlice_l165_407_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_407;
  wire       [3:0]    _zz_when_ArraySlice_l166_407_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_407_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_407_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_407_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_407;
  wire       [6:0]    _zz_when_ArraySlice_l113_407;
  wire       [6:0]    _zz_when_ArraySlice_l113_407_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_407_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_407_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_407_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_407;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_407_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_407_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_407_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_407;
  wire       [6:0]    _zz_when_ArraySlice_l118_407_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_407_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_407_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_407_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_407_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_407_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_407_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_407_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_407_8;
  wire                _zz_when_ArraySlice_l350;
  wire                _zz_when_ArraySlice_l350_1;
  wire                _zz_when_ArraySlice_l350_2;
  wire                _zz_when_ArraySlice_l350_3;
  wire                _zz_when_ArraySlice_l350_4;
  wire                _zz_when_ArraySlice_l350_5;
  wire       [5:0]    _zz_when_ArraySlice_l165_408;
  wire       [5:0]    _zz_when_ArraySlice_l165_408_1;
  wire       [2:0]    _zz_when_ArraySlice_l165_408_2;
  wire       [6:0]    _zz_when_ArraySlice_l166_408;
  wire       [6:0]    _zz_when_ArraySlice_l166_408_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_408_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_408_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_408_4;
  wire       [2:0]    _zz_when_ArraySlice_l166_408_5;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_408;
  wire       [6:0]    _zz_when_ArraySlice_l113_408;
  wire       [6:0]    _zz_when_ArraySlice_l113_408_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_408_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_408_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_408_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_408;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_408_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_408_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_408_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_408;
  wire       [6:0]    _zz_when_ArraySlice_l118_408_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_408_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_408_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_408_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_408_4;
  wire       [5:0]    _zz_when_ArraySlice_l173_408_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_408_6;
  wire       [2:0]    _zz_when_ArraySlice_l173_408_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_408_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_409;
  wire       [5:0]    _zz_when_ArraySlice_l165_409_1;
  wire       [3:0]    _zz_when_ArraySlice_l165_409_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_409;
  wire       [5:0]    _zz_when_ArraySlice_l166_409_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_409_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_409_3;
  wire       [3:0]    _zz_when_ArraySlice_l166_409_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_409;
  wire       [6:0]    _zz_when_ArraySlice_l113_409;
  wire       [6:0]    _zz_when_ArraySlice_l113_409_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_409_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_409_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_409_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_409;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_409_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_409_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_409_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_409;
  wire       [6:0]    _zz_when_ArraySlice_l118_409_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_409_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_409_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_409_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_409_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_409_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_409_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_409_7;
  wire       [3:0]    _zz_when_ArraySlice_l173_409_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_409_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_410;
  wire       [5:0]    _zz_when_ArraySlice_l165_410_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_410_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_410;
  wire       [5:0]    _zz_when_ArraySlice_l166_410_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_410_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_410_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_410_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_410;
  wire       [6:0]    _zz_when_ArraySlice_l113_410;
  wire       [6:0]    _zz_when_ArraySlice_l113_410_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_410_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_410_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_410_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_410;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_410_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_410_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_410_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_410;
  wire       [6:0]    _zz_when_ArraySlice_l118_410_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_410_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_410_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_410_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_410_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_410_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_410_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_410_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_410_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_410_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_411;
  wire       [5:0]    _zz_when_ArraySlice_l165_411_1;
  wire       [4:0]    _zz_when_ArraySlice_l165_411_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_411;
  wire       [5:0]    _zz_when_ArraySlice_l166_411_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_411_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_411_3;
  wire       [4:0]    _zz_when_ArraySlice_l166_411_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_411;
  wire       [6:0]    _zz_when_ArraySlice_l113_411;
  wire       [6:0]    _zz_when_ArraySlice_l113_411_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_411_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_411_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_411_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_411;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_411_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_411_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_411_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_411;
  wire       [6:0]    _zz_when_ArraySlice_l118_411_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_411_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_411_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_411_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_411_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_411_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_411_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_411_7;
  wire       [4:0]    _zz_when_ArraySlice_l173_411_8;
  wire       [6:0]    _zz_when_ArraySlice_l173_411_9;
  wire       [5:0]    _zz_when_ArraySlice_l165_412;
  wire       [5:0]    _zz_when_ArraySlice_l165_412_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_412;
  wire       [5:0]    _zz_when_ArraySlice_l166_412_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_412_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_412_3;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_412;
  wire       [6:0]    _zz_when_ArraySlice_l113_412;
  wire       [6:0]    _zz_when_ArraySlice_l113_412_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_412_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_412_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_412_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_412;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_412_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_412_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_412_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_412;
  wire       [6:0]    _zz_when_ArraySlice_l118_412_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_412_1;
  wire       [5:0]    _zz_when_ArraySlice_l173_412_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_412_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_412_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_412_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_412_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_412_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_412_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_413;
  wire       [5:0]    _zz_when_ArraySlice_l165_413_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_413;
  wire       [4:0]    _zz_when_ArraySlice_l166_413_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_413_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_413_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_413_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_413;
  wire       [6:0]    _zz_when_ArraySlice_l113_413;
  wire       [6:0]    _zz_when_ArraySlice_l113_413_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_413_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_413_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_413_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_413;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_413_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_413_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_413_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_413;
  wire       [6:0]    _zz_when_ArraySlice_l118_413_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_413_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_413_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_413_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_413_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_413_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_413_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_413_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_413_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_414;
  wire       [5:0]    _zz_when_ArraySlice_l165_414_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_414;
  wire       [4:0]    _zz_when_ArraySlice_l166_414_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_414_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_414_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_414_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_414;
  wire       [6:0]    _zz_when_ArraySlice_l113_414;
  wire       [6:0]    _zz_when_ArraySlice_l113_414_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_414_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_414_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_414_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_414;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_414_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_414_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_414_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_414;
  wire       [6:0]    _zz_when_ArraySlice_l118_414_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_414_1;
  wire       [4:0]    _zz_when_ArraySlice_l173_414_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_414_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_414_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_414_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_414_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_414_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_414_8;
  wire       [5:0]    _zz_when_ArraySlice_l165_415;
  wire       [5:0]    _zz_when_ArraySlice_l165_415_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_415;
  wire       [3:0]    _zz_when_ArraySlice_l166_415_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_415_2;
  wire       [5:0]    _zz_when_ArraySlice_l166_415_3;
  wire       [5:0]    _zz_when_ArraySlice_l166_415_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l112_415;
  wire       [6:0]    _zz_when_ArraySlice_l113_415;
  wire       [6:0]    _zz_when_ArraySlice_l113_415_1;
  wire       [6:0]    _zz_when_ArraySlice_l113_415_2;
  wire       [6:0]    _zz_when_ArraySlice_l113_415_3;
  wire       [6:0]    _zz_when_ArraySlice_l113_415_4;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_415;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_415_1;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_415_2;
  wire       [6:0]    _zz__zz_when_ArraySlice_l173_415_3;
  wire       [5:0]    _zz_when_ArraySlice_l118_415;
  wire       [6:0]    _zz_when_ArraySlice_l118_415_1;
  wire       [6:0]    _zz_when_ArraySlice_l173_415_1;
  wire       [3:0]    _zz_when_ArraySlice_l173_415_2;
  wire       [6:0]    _zz_when_ArraySlice_l173_415_3;
  wire       [6:0]    _zz_when_ArraySlice_l173_415_4;
  wire       [6:0]    _zz_when_ArraySlice_l173_415_5;
  wire       [5:0]    _zz_when_ArraySlice_l173_415_6;
  wire       [5:0]    _zz_when_ArraySlice_l173_415_7;
  wire       [6:0]    _zz_when_ArraySlice_l173_415_8;
  wire       [5:0]    _zz_when_ArraySlice_l189_8;
  wire       [5:0]    _zz_when_ArraySlice_l189_8_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_9;
  wire       [5:0]    _zz_when_ArraySlice_l189_9_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_10;
  wire       [5:0]    _zz_when_ArraySlice_l189_10_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_11;
  wire       [5:0]    _zz_when_ArraySlice_l189_11_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_12;
  wire       [5:0]    _zz_when_ArraySlice_l189_12_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_13;
  wire       [5:0]    _zz_when_ArraySlice_l189_13_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_14;
  wire       [5:0]    _zz_when_ArraySlice_l189_14_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_15;
  wire       [5:0]    _zz_when_ArraySlice_l189_15_1;
  wire                _zz_when_ArraySlice_l354_8;
  wire                _zz_when_ArraySlice_l354_9;
  wire                _zz_when_ArraySlice_l354_10;
  wire                _zz_when_ArraySlice_l354_11;
  wire                _zz_when_ArraySlice_l354_12;
  wire                _zz_when_ArraySlice_l354_13;
  wire                _zz_when_ArraySlice_l354_14;
  wire                _zz_when_ArraySlice_l354_15;
  wire                _zz_when_ArraySlice_l354_16;
  wire                _zz_when_ArraySlice_l354_17;
  wire                _zz_when_ArraySlice_l354_18;
  wire                _zz_when_ArraySlice_l354_19;
  wire                _zz_when_ArraySlice_l354_20;
  wire                _zz_when_ArraySlice_l354_21;
  wire                _zz_when_ArraySlice_l354_22;
  wire                _zz_when_ArraySlice_l354_23;
  wire                _zz_when_ArraySlice_l354_24;
  wire                _zz_when_ArraySlice_l354_25;
  wire       [5:0]    _zz_when_ArraySlice_l189_16;
  wire       [5:0]    _zz_when_ArraySlice_l189_16_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_17;
  wire       [5:0]    _zz_when_ArraySlice_l189_17_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_18;
  wire       [5:0]    _zz_when_ArraySlice_l189_18_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_19;
  wire       [5:0]    _zz_when_ArraySlice_l189_19_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_20;
  wire       [5:0]    _zz_when_ArraySlice_l189_20_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_21;
  wire       [5:0]    _zz_when_ArraySlice_l189_21_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_22;
  wire       [5:0]    _zz_when_ArraySlice_l189_22_1;
  wire       [5:0]    _zz_when_ArraySlice_l189_23;
  wire       [5:0]    _zz_when_ArraySlice_l189_23_1;
  wire       [31:0]   arrayDataType;
  reg        [5:0]    wReg;
  reg        [5:0]    hReg;
  reg        [2:0]    aReg;
  reg        [2:0]    bReg;
  reg                 handshakeTimes_0_willIncrement;
  reg                 handshakeTimes_0_willClear;
  reg        [12:0]   handshakeTimes_0_valueNext;
  reg        [12:0]   handshakeTimes_0_value;
  wire                handshakeTimes_0_willOverflowIfInc;
  wire                handshakeTimes_0_willOverflow;
  reg                 handshakeTimes_1_willIncrement;
  reg                 handshakeTimes_1_willClear;
  reg        [12:0]   handshakeTimes_1_valueNext;
  reg        [12:0]   handshakeTimes_1_value;
  wire                handshakeTimes_1_willOverflowIfInc;
  wire                handshakeTimes_1_willOverflow;
  reg                 handshakeTimes_2_willIncrement;
  reg                 handshakeTimes_2_willClear;
  reg        [12:0]   handshakeTimes_2_valueNext;
  reg        [12:0]   handshakeTimes_2_value;
  wire                handshakeTimes_2_willOverflowIfInc;
  wire                handshakeTimes_2_willOverflow;
  reg                 handshakeTimes_3_willIncrement;
  reg                 handshakeTimes_3_willClear;
  reg        [12:0]   handshakeTimes_3_valueNext;
  reg        [12:0]   handshakeTimes_3_value;
  wire                handshakeTimes_3_willOverflowIfInc;
  wire                handshakeTimes_3_willOverflow;
  reg                 handshakeTimes_4_willIncrement;
  reg                 handshakeTimes_4_willClear;
  reg        [12:0]   handshakeTimes_4_valueNext;
  reg        [12:0]   handshakeTimes_4_value;
  wire                handshakeTimes_4_willOverflowIfInc;
  wire                handshakeTimes_4_willOverflow;
  reg                 handshakeTimes_5_willIncrement;
  reg                 handshakeTimes_5_willClear;
  reg        [12:0]   handshakeTimes_5_valueNext;
  reg        [12:0]   handshakeTimes_5_value;
  wire                handshakeTimes_5_willOverflowIfInc;
  wire                handshakeTimes_5_willOverflow;
  reg                 handshakeTimes_6_willIncrement;
  reg                 handshakeTimes_6_willClear;
  reg        [12:0]   handshakeTimes_6_valueNext;
  reg        [12:0]   handshakeTimes_6_value;
  wire                handshakeTimes_6_willOverflowIfInc;
  wire                handshakeTimes_6_willOverflow;
  reg                 handshakeTimes_7_willIncrement;
  reg                 handshakeTimes_7_willClear;
  reg        [12:0]   handshakeTimes_7_valueNext;
  reg        [12:0]   handshakeTimes_7_value;
  wire                handshakeTimes_7_willOverflowIfInc;
  wire                handshakeTimes_7_willOverflow;
  reg        [5:0]    selectWriteFifo;
  reg        [5:0]    selectReadFifo_0;
  reg        [5:0]    selectReadFifo_1;
  reg        [5:0]    selectReadFifo_2;
  reg        [5:0]    selectReadFifo_3;
  reg        [5:0]    selectReadFifo_4;
  reg        [5:0]    selectReadFifo_5;
  reg        [5:0]    selectReadFifo_6;
  reg        [5:0]    selectReadFifo_7;
  reg                 holdReadOp_0;
  reg                 holdReadOp_1;
  reg                 holdReadOp_2;
  reg                 holdReadOp_3;
  reg                 holdReadOp_4;
  reg                 holdReadOp_5;
  reg                 holdReadOp_6;
  reg                 holdReadOp_7;
  reg                 allowPadding_0;
  reg                 allowPadding_1;
  reg                 allowPadding_2;
  reg                 allowPadding_3;
  reg                 allowPadding_4;
  reg                 allowPadding_5;
  reg                 allowPadding_6;
  reg                 allowPadding_7;
  reg                 outSliceNumb_0_willIncrement;
  reg                 outSliceNumb_0_willClear;
  reg        [6:0]    outSliceNumb_0_valueNext;
  reg        [6:0]    outSliceNumb_0_value;
  wire                outSliceNumb_0_willOverflowIfInc;
  wire                outSliceNumb_0_willOverflow;
  reg                 outSliceNumb_1_willIncrement;
  reg                 outSliceNumb_1_willClear;
  reg        [6:0]    outSliceNumb_1_valueNext;
  reg        [6:0]    outSliceNumb_1_value;
  wire                outSliceNumb_1_willOverflowIfInc;
  wire                outSliceNumb_1_willOverflow;
  reg                 outSliceNumb_2_willIncrement;
  reg                 outSliceNumb_2_willClear;
  reg        [6:0]    outSliceNumb_2_valueNext;
  reg        [6:0]    outSliceNumb_2_value;
  wire                outSliceNumb_2_willOverflowIfInc;
  wire                outSliceNumb_2_willOverflow;
  reg                 outSliceNumb_3_willIncrement;
  reg                 outSliceNumb_3_willClear;
  reg        [6:0]    outSliceNumb_3_valueNext;
  reg        [6:0]    outSliceNumb_3_value;
  wire                outSliceNumb_3_willOverflowIfInc;
  wire                outSliceNumb_3_willOverflow;
  reg                 outSliceNumb_4_willIncrement;
  reg                 outSliceNumb_4_willClear;
  reg        [6:0]    outSliceNumb_4_valueNext;
  reg        [6:0]    outSliceNumb_4_value;
  wire                outSliceNumb_4_willOverflowIfInc;
  wire                outSliceNumb_4_willOverflow;
  reg                 outSliceNumb_5_willIncrement;
  reg                 outSliceNumb_5_willClear;
  reg        [6:0]    outSliceNumb_5_valueNext;
  reg        [6:0]    outSliceNumb_5_value;
  wire                outSliceNumb_5_willOverflowIfInc;
  wire                outSliceNumb_5_willOverflow;
  reg                 outSliceNumb_6_willIncrement;
  reg                 outSliceNumb_6_willClear;
  reg        [6:0]    outSliceNumb_6_valueNext;
  reg        [6:0]    outSliceNumb_6_value;
  wire                outSliceNumb_6_willOverflowIfInc;
  wire                outSliceNumb_6_willOverflow;
  reg                 outSliceNumb_7_willIncrement;
  reg                 outSliceNumb_7_willClear;
  reg        [6:0]    outSliceNumb_7_valueNext;
  reg        [6:0]    outSliceNumb_7_value;
  wire                outSliceNumb_7_willOverflowIfInc;
  wire                outSliceNumb_7_willOverflow;
  reg                 writeAround;
  reg                 readAround_0;
  reg                 readAround_1;
  reg                 readAround_2;
  reg                 readAround_3;
  reg                 readAround_4;
  reg                 readAround_5;
  reg                 readAround_6;
  reg                 readAround_7;
  wire                arraySliceStateMachine_wantExit;
  reg                 arraySliceStateMachine_wantStart;
  wire                arraySliceStateMachine_wantKill;
  wire       [1:0]    stateIndicate;
  reg        [1:0]    arraySliceStateMachine_stateReg;
  reg        [1:0]    arraySliceStateMachine_stateNext;
  wire                when_ArraySlice_l211;
  wire                _zz_io_push_valid;
  wire       [31:0]   _zz_io_push_payload;
  wire       [63:0]   _zz_1;
  wire       [63:0]   _zz_2;
  wire                inputStreamArrayData_fire;
  wire                when_ArraySlice_l215;
  wire                when_ArraySlice_l216;
  reg                 debug_0 /* verilator public */ ;
  reg                 debug_1 /* verilator public */ ;
  reg                 debug_2 /* verilator public */ ;
  reg                 debug_3 /* verilator public */ ;
  reg                 debug_4 /* verilator public */ ;
  reg                 debug_5 /* verilator public */ ;
  reg                 debug_6 /* verilator public */ ;
  reg                 debug_7 /* verilator public */ ;
  wire                when_ArraySlice_l165;
  wire                when_ArraySlice_l166;
  reg        [6:0]    _zz_when_ArraySlice_l173;
  wire       [5:0]    _zz_when_ArraySlice_l112;
  wire                when_ArraySlice_l112;
  wire                when_ArraySlice_l113;
  wire                when_ArraySlice_l118;
  wire                when_ArraySlice_l173;
  wire                when_ArraySlice_l165_1;
  wire                when_ArraySlice_l166_1;
  reg        [6:0]    _zz_when_ArraySlice_l173_1;
  wire       [5:0]    _zz_when_ArraySlice_l112_1;
  wire                when_ArraySlice_l112_1;
  wire                when_ArraySlice_l113_1;
  wire                when_ArraySlice_l118_1;
  wire                when_ArraySlice_l173_1;
  wire                when_ArraySlice_l165_2;
  wire                when_ArraySlice_l166_2;
  reg        [6:0]    _zz_when_ArraySlice_l173_2;
  wire       [5:0]    _zz_when_ArraySlice_l112_2;
  wire                when_ArraySlice_l112_2;
  wire                when_ArraySlice_l113_2;
  wire                when_ArraySlice_l118_2;
  wire                when_ArraySlice_l173_2;
  wire                when_ArraySlice_l165_3;
  wire                when_ArraySlice_l166_3;
  reg        [6:0]    _zz_when_ArraySlice_l173_3;
  wire       [5:0]    _zz_when_ArraySlice_l112_3;
  wire                when_ArraySlice_l112_3;
  wire                when_ArraySlice_l113_3;
  wire                when_ArraySlice_l118_3;
  wire                when_ArraySlice_l173_3;
  wire                when_ArraySlice_l165_4;
  wire                when_ArraySlice_l166_4;
  reg        [6:0]    _zz_when_ArraySlice_l173_4;
  wire       [5:0]    _zz_when_ArraySlice_l112_4;
  wire                when_ArraySlice_l112_4;
  wire                when_ArraySlice_l113_4;
  wire                when_ArraySlice_l118_4;
  wire                when_ArraySlice_l173_4;
  wire                when_ArraySlice_l165_5;
  wire                when_ArraySlice_l166_5;
  reg        [6:0]    _zz_when_ArraySlice_l173_5;
  wire       [5:0]    _zz_when_ArraySlice_l112_5;
  wire                when_ArraySlice_l112_5;
  wire                when_ArraySlice_l113_5;
  wire                when_ArraySlice_l118_5;
  wire                when_ArraySlice_l173_5;
  wire                when_ArraySlice_l165_6;
  wire                when_ArraySlice_l166_6;
  reg        [6:0]    _zz_when_ArraySlice_l173_6;
  wire       [5:0]    _zz_when_ArraySlice_l112_6;
  wire                when_ArraySlice_l112_6;
  wire                when_ArraySlice_l113_6;
  wire                when_ArraySlice_l118_6;
  wire                when_ArraySlice_l173_6;
  wire                when_ArraySlice_l165_7;
  wire                when_ArraySlice_l166_7;
  reg        [6:0]    _zz_when_ArraySlice_l173_7;
  wire       [5:0]    _zz_when_ArraySlice_l112_7;
  wire                when_ArraySlice_l112_7;
  wire                when_ArraySlice_l113_7;
  wire                when_ArraySlice_l118_7;
  wire                when_ArraySlice_l173_7;
  wire                when_ArraySlice_l223;
  wire                when_ArraySlice_l229;
  wire                when_ArraySlice_l229_1;
  wire                when_ArraySlice_l229_2;
  wire                when_ArraySlice_l229_3;
  wire                when_ArraySlice_l229_4;
  wire                when_ArraySlice_l229_5;
  wire                when_ArraySlice_l229_6;
  wire                when_ArraySlice_l229_7;
  wire                when_ArraySlice_l373;
  wire                when_ArraySlice_l374;
  wire       [5:0]    _zz_outputStreamArrayData_0_valid;
  wire                _zz_io_pop_ready;
  wire       [63:0]   _zz_3;
  wire                when_ArraySlice_l379;
  wire                outputStreamArrayData_0_fire;
  wire                when_ArraySlice_l380;
  wire                when_ArraySlice_l381;
  wire                when_ArraySlice_l384;
  wire                outputStreamArrayData_0_fire_1;
  wire                when_ArraySlice_l389;
  wire                when_ArraySlice_l390;
  reg        [6:0]    _zz_when_ArraySlice_l392;
  wire       [5:0]    _zz_when_ArraySlice_l94;
  wire                when_ArraySlice_l94;
  wire                when_ArraySlice_l95;
  wire                when_ArraySlice_l99;
  wire                when_ArraySlice_l392;
  reg                 debug_0_1 /* verilator public */ ;
  reg                 debug_1_1 /* verilator public */ ;
  reg                 debug_2_1 /* verilator public */ ;
  reg                 debug_3_1 /* verilator public */ ;
  reg                 debug_4_1 /* verilator public */ ;
  reg                 debug_5_1 /* verilator public */ ;
  reg                 debug_6_1 /* verilator public */ ;
  reg                 debug_7_1 /* verilator public */ ;
  wire                when_ArraySlice_l165_8;
  wire                when_ArraySlice_l166_8;
  reg        [6:0]    _zz_when_ArraySlice_l173_8;
  wire       [5:0]    _zz_when_ArraySlice_l112_8;
  wire                when_ArraySlice_l112_8;
  wire                when_ArraySlice_l113_8;
  wire                when_ArraySlice_l118_8;
  wire                when_ArraySlice_l173_8;
  wire                when_ArraySlice_l165_9;
  wire                when_ArraySlice_l166_9;
  reg        [6:0]    _zz_when_ArraySlice_l173_9;
  wire       [5:0]    _zz_when_ArraySlice_l112_9;
  wire                when_ArraySlice_l112_9;
  wire                when_ArraySlice_l113_9;
  wire                when_ArraySlice_l118_9;
  wire                when_ArraySlice_l173_9;
  wire                when_ArraySlice_l165_10;
  wire                when_ArraySlice_l166_10;
  reg        [6:0]    _zz_when_ArraySlice_l173_10;
  wire       [5:0]    _zz_when_ArraySlice_l112_10;
  wire                when_ArraySlice_l112_10;
  wire                when_ArraySlice_l113_10;
  wire                when_ArraySlice_l118_10;
  wire                when_ArraySlice_l173_10;
  wire                when_ArraySlice_l165_11;
  wire                when_ArraySlice_l166_11;
  reg        [6:0]    _zz_when_ArraySlice_l173_11;
  wire       [5:0]    _zz_when_ArraySlice_l112_11;
  wire                when_ArraySlice_l112_11;
  wire                when_ArraySlice_l113_11;
  wire                when_ArraySlice_l118_11;
  wire                when_ArraySlice_l173_11;
  wire                when_ArraySlice_l165_12;
  wire                when_ArraySlice_l166_12;
  reg        [6:0]    _zz_when_ArraySlice_l173_12;
  wire       [5:0]    _zz_when_ArraySlice_l112_12;
  wire                when_ArraySlice_l112_12;
  wire                when_ArraySlice_l113_12;
  wire                when_ArraySlice_l118_12;
  wire                when_ArraySlice_l173_12;
  wire                when_ArraySlice_l165_13;
  wire                when_ArraySlice_l166_13;
  reg        [6:0]    _zz_when_ArraySlice_l173_13;
  wire       [5:0]    _zz_when_ArraySlice_l112_13;
  wire                when_ArraySlice_l112_13;
  wire                when_ArraySlice_l113_13;
  wire                when_ArraySlice_l118_13;
  wire                when_ArraySlice_l173_13;
  wire                when_ArraySlice_l165_14;
  wire                when_ArraySlice_l166_14;
  reg        [6:0]    _zz_when_ArraySlice_l173_14;
  wire       [5:0]    _zz_when_ArraySlice_l112_14;
  wire                when_ArraySlice_l112_14;
  wire                when_ArraySlice_l113_14;
  wire                when_ArraySlice_l118_14;
  wire                when_ArraySlice_l173_14;
  wire                when_ArraySlice_l165_15;
  wire                when_ArraySlice_l166_15;
  reg        [6:0]    _zz_when_ArraySlice_l173_15;
  wire       [5:0]    _zz_when_ArraySlice_l112_15;
  wire                when_ArraySlice_l112_15;
  wire                when_ArraySlice_l113_15;
  wire                when_ArraySlice_l118_15;
  wire                when_ArraySlice_l173_15;
  wire                when_ArraySlice_l398;
  wire                when_ArraySlice_l401;
  wire                when_ArraySlice_l405;
  wire                when_ArraySlice_l409;
  wire                outputStreamArrayData_0_fire_2;
  wire                when_ArraySlice_l410;
  reg        [6:0]    _zz_when_ArraySlice_l412;
  wire       [5:0]    _zz_when_ArraySlice_l94_1;
  wire                when_ArraySlice_l94_1;
  wire                when_ArraySlice_l95_1;
  wire                when_ArraySlice_l99_1;
  wire                when_ArraySlice_l412;
  reg                 debug_0_2 /* verilator public */ ;
  reg                 debug_1_2 /* verilator public */ ;
  reg                 debug_2_2 /* verilator public */ ;
  reg                 debug_3_2 /* verilator public */ ;
  reg                 debug_4_2 /* verilator public */ ;
  reg                 debug_5_2 /* verilator public */ ;
  reg                 debug_6_2 /* verilator public */ ;
  reg                 debug_7_2 /* verilator public */ ;
  wire                when_ArraySlice_l165_16;
  wire                when_ArraySlice_l166_16;
  reg        [6:0]    _zz_when_ArraySlice_l173_16;
  wire       [5:0]    _zz_when_ArraySlice_l112_16;
  wire                when_ArraySlice_l112_16;
  wire                when_ArraySlice_l113_16;
  wire                when_ArraySlice_l118_16;
  wire                when_ArraySlice_l173_16;
  wire                when_ArraySlice_l165_17;
  wire                when_ArraySlice_l166_17;
  reg        [6:0]    _zz_when_ArraySlice_l173_17;
  wire       [5:0]    _zz_when_ArraySlice_l112_17;
  wire                when_ArraySlice_l112_17;
  wire                when_ArraySlice_l113_17;
  wire                when_ArraySlice_l118_17;
  wire                when_ArraySlice_l173_17;
  wire                when_ArraySlice_l165_18;
  wire                when_ArraySlice_l166_18;
  reg        [6:0]    _zz_when_ArraySlice_l173_18;
  wire       [5:0]    _zz_when_ArraySlice_l112_18;
  wire                when_ArraySlice_l112_18;
  wire                when_ArraySlice_l113_18;
  wire                when_ArraySlice_l118_18;
  wire                when_ArraySlice_l173_18;
  wire                when_ArraySlice_l165_19;
  wire                when_ArraySlice_l166_19;
  reg        [6:0]    _zz_when_ArraySlice_l173_19;
  wire       [5:0]    _zz_when_ArraySlice_l112_19;
  wire                when_ArraySlice_l112_19;
  wire                when_ArraySlice_l113_19;
  wire                when_ArraySlice_l118_19;
  wire                when_ArraySlice_l173_19;
  wire                when_ArraySlice_l165_20;
  wire                when_ArraySlice_l166_20;
  reg        [6:0]    _zz_when_ArraySlice_l173_20;
  wire       [5:0]    _zz_when_ArraySlice_l112_20;
  wire                when_ArraySlice_l112_20;
  wire                when_ArraySlice_l113_20;
  wire                when_ArraySlice_l118_20;
  wire                when_ArraySlice_l173_20;
  wire                when_ArraySlice_l165_21;
  wire                when_ArraySlice_l166_21;
  reg        [6:0]    _zz_when_ArraySlice_l173_21;
  wire       [5:0]    _zz_when_ArraySlice_l112_21;
  wire                when_ArraySlice_l112_21;
  wire                when_ArraySlice_l113_21;
  wire                when_ArraySlice_l118_21;
  wire                when_ArraySlice_l173_21;
  wire                when_ArraySlice_l165_22;
  wire                when_ArraySlice_l166_22;
  reg        [6:0]    _zz_when_ArraySlice_l173_22;
  wire       [5:0]    _zz_when_ArraySlice_l112_22;
  wire                when_ArraySlice_l112_22;
  wire                when_ArraySlice_l113_22;
  wire                when_ArraySlice_l118_22;
  wire                when_ArraySlice_l173_22;
  wire                when_ArraySlice_l165_23;
  wire                when_ArraySlice_l166_23;
  reg        [6:0]    _zz_when_ArraySlice_l173_23;
  wire       [5:0]    _zz_when_ArraySlice_l112_23;
  wire                when_ArraySlice_l112_23;
  wire                when_ArraySlice_l113_23;
  wire                when_ArraySlice_l118_23;
  wire                when_ArraySlice_l173_23;
  wire                when_ArraySlice_l418;
  wire                when_ArraySlice_l421;
  wire                outputStreamArrayData_0_fire_3;
  wire                when_ArraySlice_l425;
  wire                outputStreamArrayData_0_fire_4;
  wire                when_ArraySlice_l436;
  reg        [6:0]    _zz_when_ArraySlice_l437;
  wire       [5:0]    _zz_when_ArraySlice_l94_2;
  wire                when_ArraySlice_l94_2;
  wire                when_ArraySlice_l95_2;
  wire                when_ArraySlice_l99_2;
  wire                when_ArraySlice_l437;
  reg                 debug_0_3 /* verilator public */ ;
  reg                 debug_1_3 /* verilator public */ ;
  reg                 debug_2_3 /* verilator public */ ;
  reg                 debug_3_3 /* verilator public */ ;
  reg                 debug_4_3 /* verilator public */ ;
  reg                 debug_5_3 /* verilator public */ ;
  reg                 debug_6_3 /* verilator public */ ;
  reg                 debug_7_3 /* verilator public */ ;
  wire                when_ArraySlice_l165_24;
  wire                when_ArraySlice_l166_24;
  reg        [6:0]    _zz_when_ArraySlice_l173_24;
  wire       [5:0]    _zz_when_ArraySlice_l112_24;
  wire                when_ArraySlice_l112_24;
  wire                when_ArraySlice_l113_24;
  wire                when_ArraySlice_l118_24;
  wire                when_ArraySlice_l173_24;
  wire                when_ArraySlice_l165_25;
  wire                when_ArraySlice_l166_25;
  reg        [6:0]    _zz_when_ArraySlice_l173_25;
  wire       [5:0]    _zz_when_ArraySlice_l112_25;
  wire                when_ArraySlice_l112_25;
  wire                when_ArraySlice_l113_25;
  wire                when_ArraySlice_l118_25;
  wire                when_ArraySlice_l173_25;
  wire                when_ArraySlice_l165_26;
  wire                when_ArraySlice_l166_26;
  reg        [6:0]    _zz_when_ArraySlice_l173_26;
  wire       [5:0]    _zz_when_ArraySlice_l112_26;
  wire                when_ArraySlice_l112_26;
  wire                when_ArraySlice_l113_26;
  wire                when_ArraySlice_l118_26;
  wire                when_ArraySlice_l173_26;
  wire                when_ArraySlice_l165_27;
  wire                when_ArraySlice_l166_27;
  reg        [6:0]    _zz_when_ArraySlice_l173_27;
  wire       [5:0]    _zz_when_ArraySlice_l112_27;
  wire                when_ArraySlice_l112_27;
  wire                when_ArraySlice_l113_27;
  wire                when_ArraySlice_l118_27;
  wire                when_ArraySlice_l173_27;
  wire                when_ArraySlice_l165_28;
  wire                when_ArraySlice_l166_28;
  reg        [6:0]    _zz_when_ArraySlice_l173_28;
  wire       [5:0]    _zz_when_ArraySlice_l112_28;
  wire                when_ArraySlice_l112_28;
  wire                when_ArraySlice_l113_28;
  wire                when_ArraySlice_l118_28;
  wire                when_ArraySlice_l173_28;
  wire                when_ArraySlice_l165_29;
  wire                when_ArraySlice_l166_29;
  reg        [6:0]    _zz_when_ArraySlice_l173_29;
  wire       [5:0]    _zz_when_ArraySlice_l112_29;
  wire                when_ArraySlice_l112_29;
  wire                when_ArraySlice_l113_29;
  wire                when_ArraySlice_l118_29;
  wire                when_ArraySlice_l173_29;
  wire                when_ArraySlice_l165_30;
  wire                when_ArraySlice_l166_30;
  reg        [6:0]    _zz_when_ArraySlice_l173_30;
  wire       [5:0]    _zz_when_ArraySlice_l112_30;
  wire                when_ArraySlice_l112_30;
  wire                when_ArraySlice_l113_30;
  wire                when_ArraySlice_l118_30;
  wire                when_ArraySlice_l173_30;
  wire                when_ArraySlice_l165_31;
  wire                when_ArraySlice_l166_31;
  reg        [6:0]    _zz_when_ArraySlice_l173_31;
  wire       [5:0]    _zz_when_ArraySlice_l112_31;
  wire                when_ArraySlice_l112_31;
  wire                when_ArraySlice_l113_31;
  wire                when_ArraySlice_l118_31;
  wire                when_ArraySlice_l173_31;
  wire                when_ArraySlice_l444;
  wire                outputStreamArrayData_0_fire_5;
  wire                when_ArraySlice_l448;
  wire                when_ArraySlice_l434;
  wire                outputStreamArrayData_0_fire_6;
  wire                when_ArraySlice_l455;
  wire                when_ArraySlice_l373_1;
  wire                when_ArraySlice_l374_1;
  wire       [5:0]    _zz_outputStreamArrayData_1_valid;
  wire                _zz_io_pop_ready_1;
  wire       [63:0]   _zz_4;
  wire                when_ArraySlice_l379_1;
  wire                outputStreamArrayData_1_fire;
  wire                when_ArraySlice_l380_1;
  wire                when_ArraySlice_l381_1;
  wire                when_ArraySlice_l384_1;
  wire                outputStreamArrayData_1_fire_1;
  wire                when_ArraySlice_l389_1;
  wire                when_ArraySlice_l390_1;
  reg        [6:0]    _zz_when_ArraySlice_l392_1;
  wire       [5:0]    _zz_when_ArraySlice_l94_3;
  wire                when_ArraySlice_l94_3;
  wire                when_ArraySlice_l95_3;
  wire                when_ArraySlice_l99_3;
  wire                when_ArraySlice_l392_1;
  reg                 debug_0_4 /* verilator public */ ;
  reg                 debug_1_4 /* verilator public */ ;
  reg                 debug_2_4 /* verilator public */ ;
  reg                 debug_3_4 /* verilator public */ ;
  reg                 debug_4_4 /* verilator public */ ;
  reg                 debug_5_4 /* verilator public */ ;
  reg                 debug_6_4 /* verilator public */ ;
  reg                 debug_7_4 /* verilator public */ ;
  wire                when_ArraySlice_l165_32;
  wire                when_ArraySlice_l166_32;
  reg        [6:0]    _zz_when_ArraySlice_l173_32;
  wire       [5:0]    _zz_when_ArraySlice_l112_32;
  wire                when_ArraySlice_l112_32;
  wire                when_ArraySlice_l113_32;
  wire                when_ArraySlice_l118_32;
  wire                when_ArraySlice_l173_32;
  wire                when_ArraySlice_l165_33;
  wire                when_ArraySlice_l166_33;
  reg        [6:0]    _zz_when_ArraySlice_l173_33;
  wire       [5:0]    _zz_when_ArraySlice_l112_33;
  wire                when_ArraySlice_l112_33;
  wire                when_ArraySlice_l113_33;
  wire                when_ArraySlice_l118_33;
  wire                when_ArraySlice_l173_33;
  wire                when_ArraySlice_l165_34;
  wire                when_ArraySlice_l166_34;
  reg        [6:0]    _zz_when_ArraySlice_l173_34;
  wire       [5:0]    _zz_when_ArraySlice_l112_34;
  wire                when_ArraySlice_l112_34;
  wire                when_ArraySlice_l113_34;
  wire                when_ArraySlice_l118_34;
  wire                when_ArraySlice_l173_34;
  wire                when_ArraySlice_l165_35;
  wire                when_ArraySlice_l166_35;
  reg        [6:0]    _zz_when_ArraySlice_l173_35;
  wire       [5:0]    _zz_when_ArraySlice_l112_35;
  wire                when_ArraySlice_l112_35;
  wire                when_ArraySlice_l113_35;
  wire                when_ArraySlice_l118_35;
  wire                when_ArraySlice_l173_35;
  wire                when_ArraySlice_l165_36;
  wire                when_ArraySlice_l166_36;
  reg        [6:0]    _zz_when_ArraySlice_l173_36;
  wire       [5:0]    _zz_when_ArraySlice_l112_36;
  wire                when_ArraySlice_l112_36;
  wire                when_ArraySlice_l113_36;
  wire                when_ArraySlice_l118_36;
  wire                when_ArraySlice_l173_36;
  wire                when_ArraySlice_l165_37;
  wire                when_ArraySlice_l166_37;
  reg        [6:0]    _zz_when_ArraySlice_l173_37;
  wire       [5:0]    _zz_when_ArraySlice_l112_37;
  wire                when_ArraySlice_l112_37;
  wire                when_ArraySlice_l113_37;
  wire                when_ArraySlice_l118_37;
  wire                when_ArraySlice_l173_37;
  wire                when_ArraySlice_l165_38;
  wire                when_ArraySlice_l166_38;
  reg        [6:0]    _zz_when_ArraySlice_l173_38;
  wire       [5:0]    _zz_when_ArraySlice_l112_38;
  wire                when_ArraySlice_l112_38;
  wire                when_ArraySlice_l113_38;
  wire                when_ArraySlice_l118_38;
  wire                when_ArraySlice_l173_38;
  wire                when_ArraySlice_l165_39;
  wire                when_ArraySlice_l166_39;
  reg        [6:0]    _zz_when_ArraySlice_l173_39;
  wire       [5:0]    _zz_when_ArraySlice_l112_39;
  wire                when_ArraySlice_l112_39;
  wire                when_ArraySlice_l113_39;
  wire                when_ArraySlice_l118_39;
  wire                when_ArraySlice_l173_39;
  wire                when_ArraySlice_l398_1;
  wire                when_ArraySlice_l401_1;
  wire                when_ArraySlice_l405_1;
  wire                when_ArraySlice_l409_1;
  wire                outputStreamArrayData_1_fire_2;
  wire                when_ArraySlice_l410_1;
  reg        [6:0]    _zz_when_ArraySlice_l412_1;
  wire       [5:0]    _zz_when_ArraySlice_l94_4;
  wire                when_ArraySlice_l94_4;
  wire                when_ArraySlice_l95_4;
  wire                when_ArraySlice_l99_4;
  wire                when_ArraySlice_l412_1;
  reg                 debug_0_5 /* verilator public */ ;
  reg                 debug_1_5 /* verilator public */ ;
  reg                 debug_2_5 /* verilator public */ ;
  reg                 debug_3_5 /* verilator public */ ;
  reg                 debug_4_5 /* verilator public */ ;
  reg                 debug_5_5 /* verilator public */ ;
  reg                 debug_6_5 /* verilator public */ ;
  reg                 debug_7_5 /* verilator public */ ;
  wire                when_ArraySlice_l165_40;
  wire                when_ArraySlice_l166_40;
  reg        [6:0]    _zz_when_ArraySlice_l173_40;
  wire       [5:0]    _zz_when_ArraySlice_l112_40;
  wire                when_ArraySlice_l112_40;
  wire                when_ArraySlice_l113_40;
  wire                when_ArraySlice_l118_40;
  wire                when_ArraySlice_l173_40;
  wire                when_ArraySlice_l165_41;
  wire                when_ArraySlice_l166_41;
  reg        [6:0]    _zz_when_ArraySlice_l173_41;
  wire       [5:0]    _zz_when_ArraySlice_l112_41;
  wire                when_ArraySlice_l112_41;
  wire                when_ArraySlice_l113_41;
  wire                when_ArraySlice_l118_41;
  wire                when_ArraySlice_l173_41;
  wire                when_ArraySlice_l165_42;
  wire                when_ArraySlice_l166_42;
  reg        [6:0]    _zz_when_ArraySlice_l173_42;
  wire       [5:0]    _zz_when_ArraySlice_l112_42;
  wire                when_ArraySlice_l112_42;
  wire                when_ArraySlice_l113_42;
  wire                when_ArraySlice_l118_42;
  wire                when_ArraySlice_l173_42;
  wire                when_ArraySlice_l165_43;
  wire                when_ArraySlice_l166_43;
  reg        [6:0]    _zz_when_ArraySlice_l173_43;
  wire       [5:0]    _zz_when_ArraySlice_l112_43;
  wire                when_ArraySlice_l112_43;
  wire                when_ArraySlice_l113_43;
  wire                when_ArraySlice_l118_43;
  wire                when_ArraySlice_l173_43;
  wire                when_ArraySlice_l165_44;
  wire                when_ArraySlice_l166_44;
  reg        [6:0]    _zz_when_ArraySlice_l173_44;
  wire       [5:0]    _zz_when_ArraySlice_l112_44;
  wire                when_ArraySlice_l112_44;
  wire                when_ArraySlice_l113_44;
  wire                when_ArraySlice_l118_44;
  wire                when_ArraySlice_l173_44;
  wire                when_ArraySlice_l165_45;
  wire                when_ArraySlice_l166_45;
  reg        [6:0]    _zz_when_ArraySlice_l173_45;
  wire       [5:0]    _zz_when_ArraySlice_l112_45;
  wire                when_ArraySlice_l112_45;
  wire                when_ArraySlice_l113_45;
  wire                when_ArraySlice_l118_45;
  wire                when_ArraySlice_l173_45;
  wire                when_ArraySlice_l165_46;
  wire                when_ArraySlice_l166_46;
  reg        [6:0]    _zz_when_ArraySlice_l173_46;
  wire       [5:0]    _zz_when_ArraySlice_l112_46;
  wire                when_ArraySlice_l112_46;
  wire                when_ArraySlice_l113_46;
  wire                when_ArraySlice_l118_46;
  wire                when_ArraySlice_l173_46;
  wire                when_ArraySlice_l165_47;
  wire                when_ArraySlice_l166_47;
  reg        [6:0]    _zz_when_ArraySlice_l173_47;
  wire       [5:0]    _zz_when_ArraySlice_l112_47;
  wire                when_ArraySlice_l112_47;
  wire                when_ArraySlice_l113_47;
  wire                when_ArraySlice_l118_47;
  wire                when_ArraySlice_l173_47;
  wire                when_ArraySlice_l418_1;
  wire                when_ArraySlice_l421_1;
  wire                outputStreamArrayData_1_fire_3;
  wire                when_ArraySlice_l425_1;
  wire                outputStreamArrayData_1_fire_4;
  wire                when_ArraySlice_l436_1;
  reg        [6:0]    _zz_when_ArraySlice_l437_1;
  wire       [5:0]    _zz_when_ArraySlice_l94_5;
  wire                when_ArraySlice_l94_5;
  wire                when_ArraySlice_l95_5;
  wire                when_ArraySlice_l99_5;
  wire                when_ArraySlice_l437_1;
  reg                 debug_0_6 /* verilator public */ ;
  reg                 debug_1_6 /* verilator public */ ;
  reg                 debug_2_6 /* verilator public */ ;
  reg                 debug_3_6 /* verilator public */ ;
  reg                 debug_4_6 /* verilator public */ ;
  reg                 debug_5_6 /* verilator public */ ;
  reg                 debug_6_6 /* verilator public */ ;
  reg                 debug_7_6 /* verilator public */ ;
  wire                when_ArraySlice_l165_48;
  wire                when_ArraySlice_l166_48;
  reg        [6:0]    _zz_when_ArraySlice_l173_48;
  wire       [5:0]    _zz_when_ArraySlice_l112_48;
  wire                when_ArraySlice_l112_48;
  wire                when_ArraySlice_l113_48;
  wire                when_ArraySlice_l118_48;
  wire                when_ArraySlice_l173_48;
  wire                when_ArraySlice_l165_49;
  wire                when_ArraySlice_l166_49;
  reg        [6:0]    _zz_when_ArraySlice_l173_49;
  wire       [5:0]    _zz_when_ArraySlice_l112_49;
  wire                when_ArraySlice_l112_49;
  wire                when_ArraySlice_l113_49;
  wire                when_ArraySlice_l118_49;
  wire                when_ArraySlice_l173_49;
  wire                when_ArraySlice_l165_50;
  wire                when_ArraySlice_l166_50;
  reg        [6:0]    _zz_when_ArraySlice_l173_50;
  wire       [5:0]    _zz_when_ArraySlice_l112_50;
  wire                when_ArraySlice_l112_50;
  wire                when_ArraySlice_l113_50;
  wire                when_ArraySlice_l118_50;
  wire                when_ArraySlice_l173_50;
  wire                when_ArraySlice_l165_51;
  wire                when_ArraySlice_l166_51;
  reg        [6:0]    _zz_when_ArraySlice_l173_51;
  wire       [5:0]    _zz_when_ArraySlice_l112_51;
  wire                when_ArraySlice_l112_51;
  wire                when_ArraySlice_l113_51;
  wire                when_ArraySlice_l118_51;
  wire                when_ArraySlice_l173_51;
  wire                when_ArraySlice_l165_52;
  wire                when_ArraySlice_l166_52;
  reg        [6:0]    _zz_when_ArraySlice_l173_52;
  wire       [5:0]    _zz_when_ArraySlice_l112_52;
  wire                when_ArraySlice_l112_52;
  wire                when_ArraySlice_l113_52;
  wire                when_ArraySlice_l118_52;
  wire                when_ArraySlice_l173_52;
  wire                when_ArraySlice_l165_53;
  wire                when_ArraySlice_l166_53;
  reg        [6:0]    _zz_when_ArraySlice_l173_53;
  wire       [5:0]    _zz_when_ArraySlice_l112_53;
  wire                when_ArraySlice_l112_53;
  wire                when_ArraySlice_l113_53;
  wire                when_ArraySlice_l118_53;
  wire                when_ArraySlice_l173_53;
  wire                when_ArraySlice_l165_54;
  wire                when_ArraySlice_l166_54;
  reg        [6:0]    _zz_when_ArraySlice_l173_54;
  wire       [5:0]    _zz_when_ArraySlice_l112_54;
  wire                when_ArraySlice_l112_54;
  wire                when_ArraySlice_l113_54;
  wire                when_ArraySlice_l118_54;
  wire                when_ArraySlice_l173_54;
  wire                when_ArraySlice_l165_55;
  wire                when_ArraySlice_l166_55;
  reg        [6:0]    _zz_when_ArraySlice_l173_55;
  wire       [5:0]    _zz_when_ArraySlice_l112_55;
  wire                when_ArraySlice_l112_55;
  wire                when_ArraySlice_l113_55;
  wire                when_ArraySlice_l118_55;
  wire                when_ArraySlice_l173_55;
  wire                when_ArraySlice_l444_1;
  wire                outputStreamArrayData_1_fire_5;
  wire                when_ArraySlice_l448_1;
  wire                when_ArraySlice_l434_1;
  wire                outputStreamArrayData_1_fire_6;
  wire                when_ArraySlice_l455_1;
  wire                when_ArraySlice_l373_2;
  wire                when_ArraySlice_l374_2;
  wire       [5:0]    _zz_outputStreamArrayData_2_valid;
  wire                _zz_io_pop_ready_2;
  wire       [63:0]   _zz_5;
  wire                when_ArraySlice_l379_2;
  wire                outputStreamArrayData_2_fire;
  wire                when_ArraySlice_l380_2;
  wire                when_ArraySlice_l381_2;
  wire                when_ArraySlice_l384_2;
  wire                outputStreamArrayData_2_fire_1;
  wire                when_ArraySlice_l389_2;
  wire                when_ArraySlice_l390_2;
  reg        [6:0]    _zz_when_ArraySlice_l392_2;
  wire       [5:0]    _zz_when_ArraySlice_l94_6;
  wire                when_ArraySlice_l94_6;
  wire                when_ArraySlice_l95_6;
  wire                when_ArraySlice_l99_6;
  wire                when_ArraySlice_l392_2;
  reg                 debug_0_7 /* verilator public */ ;
  reg                 debug_1_7 /* verilator public */ ;
  reg                 debug_2_7 /* verilator public */ ;
  reg                 debug_3_7 /* verilator public */ ;
  reg                 debug_4_7 /* verilator public */ ;
  reg                 debug_5_7 /* verilator public */ ;
  reg                 debug_6_7 /* verilator public */ ;
  reg                 debug_7_7 /* verilator public */ ;
  wire                when_ArraySlice_l165_56;
  wire                when_ArraySlice_l166_56;
  reg        [6:0]    _zz_when_ArraySlice_l173_56;
  wire       [5:0]    _zz_when_ArraySlice_l112_56;
  wire                when_ArraySlice_l112_56;
  wire                when_ArraySlice_l113_56;
  wire                when_ArraySlice_l118_56;
  wire                when_ArraySlice_l173_56;
  wire                when_ArraySlice_l165_57;
  wire                when_ArraySlice_l166_57;
  reg        [6:0]    _zz_when_ArraySlice_l173_57;
  wire       [5:0]    _zz_when_ArraySlice_l112_57;
  wire                when_ArraySlice_l112_57;
  wire                when_ArraySlice_l113_57;
  wire                when_ArraySlice_l118_57;
  wire                when_ArraySlice_l173_57;
  wire                when_ArraySlice_l165_58;
  wire                when_ArraySlice_l166_58;
  reg        [6:0]    _zz_when_ArraySlice_l173_58;
  wire       [5:0]    _zz_when_ArraySlice_l112_58;
  wire                when_ArraySlice_l112_58;
  wire                when_ArraySlice_l113_58;
  wire                when_ArraySlice_l118_58;
  wire                when_ArraySlice_l173_58;
  wire                when_ArraySlice_l165_59;
  wire                when_ArraySlice_l166_59;
  reg        [6:0]    _zz_when_ArraySlice_l173_59;
  wire       [5:0]    _zz_when_ArraySlice_l112_59;
  wire                when_ArraySlice_l112_59;
  wire                when_ArraySlice_l113_59;
  wire                when_ArraySlice_l118_59;
  wire                when_ArraySlice_l173_59;
  wire                when_ArraySlice_l165_60;
  wire                when_ArraySlice_l166_60;
  reg        [6:0]    _zz_when_ArraySlice_l173_60;
  wire       [5:0]    _zz_when_ArraySlice_l112_60;
  wire                when_ArraySlice_l112_60;
  wire                when_ArraySlice_l113_60;
  wire                when_ArraySlice_l118_60;
  wire                when_ArraySlice_l173_60;
  wire                when_ArraySlice_l165_61;
  wire                when_ArraySlice_l166_61;
  reg        [6:0]    _zz_when_ArraySlice_l173_61;
  wire       [5:0]    _zz_when_ArraySlice_l112_61;
  wire                when_ArraySlice_l112_61;
  wire                when_ArraySlice_l113_61;
  wire                when_ArraySlice_l118_61;
  wire                when_ArraySlice_l173_61;
  wire                when_ArraySlice_l165_62;
  wire                when_ArraySlice_l166_62;
  reg        [6:0]    _zz_when_ArraySlice_l173_62;
  wire       [5:0]    _zz_when_ArraySlice_l112_62;
  wire                when_ArraySlice_l112_62;
  wire                when_ArraySlice_l113_62;
  wire                when_ArraySlice_l118_62;
  wire                when_ArraySlice_l173_62;
  wire                when_ArraySlice_l165_63;
  wire                when_ArraySlice_l166_63;
  reg        [6:0]    _zz_when_ArraySlice_l173_63;
  wire       [5:0]    _zz_when_ArraySlice_l112_63;
  wire                when_ArraySlice_l112_63;
  wire                when_ArraySlice_l113_63;
  wire                when_ArraySlice_l118_63;
  wire                when_ArraySlice_l173_63;
  wire                when_ArraySlice_l398_2;
  wire                when_ArraySlice_l401_2;
  wire                when_ArraySlice_l405_2;
  wire                when_ArraySlice_l409_2;
  wire                outputStreamArrayData_2_fire_2;
  wire                when_ArraySlice_l410_2;
  reg        [6:0]    _zz_when_ArraySlice_l412_2;
  wire       [5:0]    _zz_when_ArraySlice_l94_7;
  wire                when_ArraySlice_l94_7;
  wire                when_ArraySlice_l95_7;
  wire                when_ArraySlice_l99_7;
  wire                when_ArraySlice_l412_2;
  reg                 debug_0_8 /* verilator public */ ;
  reg                 debug_1_8 /* verilator public */ ;
  reg                 debug_2_8 /* verilator public */ ;
  reg                 debug_3_8 /* verilator public */ ;
  reg                 debug_4_8 /* verilator public */ ;
  reg                 debug_5_8 /* verilator public */ ;
  reg                 debug_6_8 /* verilator public */ ;
  reg                 debug_7_8 /* verilator public */ ;
  wire                when_ArraySlice_l165_64;
  wire                when_ArraySlice_l166_64;
  reg        [6:0]    _zz_when_ArraySlice_l173_64;
  wire       [5:0]    _zz_when_ArraySlice_l112_64;
  wire                when_ArraySlice_l112_64;
  wire                when_ArraySlice_l113_64;
  wire                when_ArraySlice_l118_64;
  wire                when_ArraySlice_l173_64;
  wire                when_ArraySlice_l165_65;
  wire                when_ArraySlice_l166_65;
  reg        [6:0]    _zz_when_ArraySlice_l173_65;
  wire       [5:0]    _zz_when_ArraySlice_l112_65;
  wire                when_ArraySlice_l112_65;
  wire                when_ArraySlice_l113_65;
  wire                when_ArraySlice_l118_65;
  wire                when_ArraySlice_l173_65;
  wire                when_ArraySlice_l165_66;
  wire                when_ArraySlice_l166_66;
  reg        [6:0]    _zz_when_ArraySlice_l173_66;
  wire       [5:0]    _zz_when_ArraySlice_l112_66;
  wire                when_ArraySlice_l112_66;
  wire                when_ArraySlice_l113_66;
  wire                when_ArraySlice_l118_66;
  wire                when_ArraySlice_l173_66;
  wire                when_ArraySlice_l165_67;
  wire                when_ArraySlice_l166_67;
  reg        [6:0]    _zz_when_ArraySlice_l173_67;
  wire       [5:0]    _zz_when_ArraySlice_l112_67;
  wire                when_ArraySlice_l112_67;
  wire                when_ArraySlice_l113_67;
  wire                when_ArraySlice_l118_67;
  wire                when_ArraySlice_l173_67;
  wire                when_ArraySlice_l165_68;
  wire                when_ArraySlice_l166_68;
  reg        [6:0]    _zz_when_ArraySlice_l173_68;
  wire       [5:0]    _zz_when_ArraySlice_l112_68;
  wire                when_ArraySlice_l112_68;
  wire                when_ArraySlice_l113_68;
  wire                when_ArraySlice_l118_68;
  wire                when_ArraySlice_l173_68;
  wire                when_ArraySlice_l165_69;
  wire                when_ArraySlice_l166_69;
  reg        [6:0]    _zz_when_ArraySlice_l173_69;
  wire       [5:0]    _zz_when_ArraySlice_l112_69;
  wire                when_ArraySlice_l112_69;
  wire                when_ArraySlice_l113_69;
  wire                when_ArraySlice_l118_69;
  wire                when_ArraySlice_l173_69;
  wire                when_ArraySlice_l165_70;
  wire                when_ArraySlice_l166_70;
  reg        [6:0]    _zz_when_ArraySlice_l173_70;
  wire       [5:0]    _zz_when_ArraySlice_l112_70;
  wire                when_ArraySlice_l112_70;
  wire                when_ArraySlice_l113_70;
  wire                when_ArraySlice_l118_70;
  wire                when_ArraySlice_l173_70;
  wire                when_ArraySlice_l165_71;
  wire                when_ArraySlice_l166_71;
  reg        [6:0]    _zz_when_ArraySlice_l173_71;
  wire       [5:0]    _zz_when_ArraySlice_l112_71;
  wire                when_ArraySlice_l112_71;
  wire                when_ArraySlice_l113_71;
  wire                when_ArraySlice_l118_71;
  wire                when_ArraySlice_l173_71;
  wire                when_ArraySlice_l418_2;
  wire                when_ArraySlice_l421_2;
  wire                outputStreamArrayData_2_fire_3;
  wire                when_ArraySlice_l425_2;
  wire                outputStreamArrayData_2_fire_4;
  wire                when_ArraySlice_l436_2;
  reg        [6:0]    _zz_when_ArraySlice_l437_2;
  wire       [5:0]    _zz_when_ArraySlice_l94_8;
  wire                when_ArraySlice_l94_8;
  wire                when_ArraySlice_l95_8;
  wire                when_ArraySlice_l99_8;
  wire                when_ArraySlice_l437_2;
  reg                 debug_0_9 /* verilator public */ ;
  reg                 debug_1_9 /* verilator public */ ;
  reg                 debug_2_9 /* verilator public */ ;
  reg                 debug_3_9 /* verilator public */ ;
  reg                 debug_4_9 /* verilator public */ ;
  reg                 debug_5_9 /* verilator public */ ;
  reg                 debug_6_9 /* verilator public */ ;
  reg                 debug_7_9 /* verilator public */ ;
  wire                when_ArraySlice_l165_72;
  wire                when_ArraySlice_l166_72;
  reg        [6:0]    _zz_when_ArraySlice_l173_72;
  wire       [5:0]    _zz_when_ArraySlice_l112_72;
  wire                when_ArraySlice_l112_72;
  wire                when_ArraySlice_l113_72;
  wire                when_ArraySlice_l118_72;
  wire                when_ArraySlice_l173_72;
  wire                when_ArraySlice_l165_73;
  wire                when_ArraySlice_l166_73;
  reg        [6:0]    _zz_when_ArraySlice_l173_73;
  wire       [5:0]    _zz_when_ArraySlice_l112_73;
  wire                when_ArraySlice_l112_73;
  wire                when_ArraySlice_l113_73;
  wire                when_ArraySlice_l118_73;
  wire                when_ArraySlice_l173_73;
  wire                when_ArraySlice_l165_74;
  wire                when_ArraySlice_l166_74;
  reg        [6:0]    _zz_when_ArraySlice_l173_74;
  wire       [5:0]    _zz_when_ArraySlice_l112_74;
  wire                when_ArraySlice_l112_74;
  wire                when_ArraySlice_l113_74;
  wire                when_ArraySlice_l118_74;
  wire                when_ArraySlice_l173_74;
  wire                when_ArraySlice_l165_75;
  wire                when_ArraySlice_l166_75;
  reg        [6:0]    _zz_when_ArraySlice_l173_75;
  wire       [5:0]    _zz_when_ArraySlice_l112_75;
  wire                when_ArraySlice_l112_75;
  wire                when_ArraySlice_l113_75;
  wire                when_ArraySlice_l118_75;
  wire                when_ArraySlice_l173_75;
  wire                when_ArraySlice_l165_76;
  wire                when_ArraySlice_l166_76;
  reg        [6:0]    _zz_when_ArraySlice_l173_76;
  wire       [5:0]    _zz_when_ArraySlice_l112_76;
  wire                when_ArraySlice_l112_76;
  wire                when_ArraySlice_l113_76;
  wire                when_ArraySlice_l118_76;
  wire                when_ArraySlice_l173_76;
  wire                when_ArraySlice_l165_77;
  wire                when_ArraySlice_l166_77;
  reg        [6:0]    _zz_when_ArraySlice_l173_77;
  wire       [5:0]    _zz_when_ArraySlice_l112_77;
  wire                when_ArraySlice_l112_77;
  wire                when_ArraySlice_l113_77;
  wire                when_ArraySlice_l118_77;
  wire                when_ArraySlice_l173_77;
  wire                when_ArraySlice_l165_78;
  wire                when_ArraySlice_l166_78;
  reg        [6:0]    _zz_when_ArraySlice_l173_78;
  wire       [5:0]    _zz_when_ArraySlice_l112_78;
  wire                when_ArraySlice_l112_78;
  wire                when_ArraySlice_l113_78;
  wire                when_ArraySlice_l118_78;
  wire                when_ArraySlice_l173_78;
  wire                when_ArraySlice_l165_79;
  wire                when_ArraySlice_l166_79;
  reg        [6:0]    _zz_when_ArraySlice_l173_79;
  wire       [5:0]    _zz_when_ArraySlice_l112_79;
  wire                when_ArraySlice_l112_79;
  wire                when_ArraySlice_l113_79;
  wire                when_ArraySlice_l118_79;
  wire                when_ArraySlice_l173_79;
  wire                when_ArraySlice_l444_2;
  wire                outputStreamArrayData_2_fire_5;
  wire                when_ArraySlice_l448_2;
  wire                when_ArraySlice_l434_2;
  wire                outputStreamArrayData_2_fire_6;
  wire                when_ArraySlice_l455_2;
  wire                when_ArraySlice_l373_3;
  wire                when_ArraySlice_l374_3;
  wire       [5:0]    _zz_outputStreamArrayData_3_valid;
  wire                _zz_io_pop_ready_3;
  wire       [63:0]   _zz_6;
  wire                when_ArraySlice_l379_3;
  wire                outputStreamArrayData_3_fire;
  wire                when_ArraySlice_l380_3;
  wire                when_ArraySlice_l381_3;
  wire                when_ArraySlice_l384_3;
  wire                outputStreamArrayData_3_fire_1;
  wire                when_ArraySlice_l389_3;
  wire                when_ArraySlice_l390_3;
  reg        [6:0]    _zz_when_ArraySlice_l392_3;
  wire       [5:0]    _zz_when_ArraySlice_l94_9;
  wire                when_ArraySlice_l94_9;
  wire                when_ArraySlice_l95_9;
  wire                when_ArraySlice_l99_9;
  wire                when_ArraySlice_l392_3;
  reg                 debug_0_10 /* verilator public */ ;
  reg                 debug_1_10 /* verilator public */ ;
  reg                 debug_2_10 /* verilator public */ ;
  reg                 debug_3_10 /* verilator public */ ;
  reg                 debug_4_10 /* verilator public */ ;
  reg                 debug_5_10 /* verilator public */ ;
  reg                 debug_6_10 /* verilator public */ ;
  reg                 debug_7_10 /* verilator public */ ;
  wire                when_ArraySlice_l165_80;
  wire                when_ArraySlice_l166_80;
  reg        [6:0]    _zz_when_ArraySlice_l173_80;
  wire       [5:0]    _zz_when_ArraySlice_l112_80;
  wire                when_ArraySlice_l112_80;
  wire                when_ArraySlice_l113_80;
  wire                when_ArraySlice_l118_80;
  wire                when_ArraySlice_l173_80;
  wire                when_ArraySlice_l165_81;
  wire                when_ArraySlice_l166_81;
  reg        [6:0]    _zz_when_ArraySlice_l173_81;
  wire       [5:0]    _zz_when_ArraySlice_l112_81;
  wire                when_ArraySlice_l112_81;
  wire                when_ArraySlice_l113_81;
  wire                when_ArraySlice_l118_81;
  wire                when_ArraySlice_l173_81;
  wire                when_ArraySlice_l165_82;
  wire                when_ArraySlice_l166_82;
  reg        [6:0]    _zz_when_ArraySlice_l173_82;
  wire       [5:0]    _zz_when_ArraySlice_l112_82;
  wire                when_ArraySlice_l112_82;
  wire                when_ArraySlice_l113_82;
  wire                when_ArraySlice_l118_82;
  wire                when_ArraySlice_l173_82;
  wire                when_ArraySlice_l165_83;
  wire                when_ArraySlice_l166_83;
  reg        [6:0]    _zz_when_ArraySlice_l173_83;
  wire       [5:0]    _zz_when_ArraySlice_l112_83;
  wire                when_ArraySlice_l112_83;
  wire                when_ArraySlice_l113_83;
  wire                when_ArraySlice_l118_83;
  wire                when_ArraySlice_l173_83;
  wire                when_ArraySlice_l165_84;
  wire                when_ArraySlice_l166_84;
  reg        [6:0]    _zz_when_ArraySlice_l173_84;
  wire       [5:0]    _zz_when_ArraySlice_l112_84;
  wire                when_ArraySlice_l112_84;
  wire                when_ArraySlice_l113_84;
  wire                when_ArraySlice_l118_84;
  wire                when_ArraySlice_l173_84;
  wire                when_ArraySlice_l165_85;
  wire                when_ArraySlice_l166_85;
  reg        [6:0]    _zz_when_ArraySlice_l173_85;
  wire       [5:0]    _zz_when_ArraySlice_l112_85;
  wire                when_ArraySlice_l112_85;
  wire                when_ArraySlice_l113_85;
  wire                when_ArraySlice_l118_85;
  wire                when_ArraySlice_l173_85;
  wire                when_ArraySlice_l165_86;
  wire                when_ArraySlice_l166_86;
  reg        [6:0]    _zz_when_ArraySlice_l173_86;
  wire       [5:0]    _zz_when_ArraySlice_l112_86;
  wire                when_ArraySlice_l112_86;
  wire                when_ArraySlice_l113_86;
  wire                when_ArraySlice_l118_86;
  wire                when_ArraySlice_l173_86;
  wire                when_ArraySlice_l165_87;
  wire                when_ArraySlice_l166_87;
  reg        [6:0]    _zz_when_ArraySlice_l173_87;
  wire       [5:0]    _zz_when_ArraySlice_l112_87;
  wire                when_ArraySlice_l112_87;
  wire                when_ArraySlice_l113_87;
  wire                when_ArraySlice_l118_87;
  wire                when_ArraySlice_l173_87;
  wire                when_ArraySlice_l398_3;
  wire                when_ArraySlice_l401_3;
  wire                when_ArraySlice_l405_3;
  wire                when_ArraySlice_l409_3;
  wire                outputStreamArrayData_3_fire_2;
  wire                when_ArraySlice_l410_3;
  reg        [6:0]    _zz_when_ArraySlice_l412_3;
  wire       [5:0]    _zz_when_ArraySlice_l94_10;
  wire                when_ArraySlice_l94_10;
  wire                when_ArraySlice_l95_10;
  wire                when_ArraySlice_l99_10;
  wire                when_ArraySlice_l412_3;
  reg                 debug_0_11 /* verilator public */ ;
  reg                 debug_1_11 /* verilator public */ ;
  reg                 debug_2_11 /* verilator public */ ;
  reg                 debug_3_11 /* verilator public */ ;
  reg                 debug_4_11 /* verilator public */ ;
  reg                 debug_5_11 /* verilator public */ ;
  reg                 debug_6_11 /* verilator public */ ;
  reg                 debug_7_11 /* verilator public */ ;
  wire                when_ArraySlice_l165_88;
  wire                when_ArraySlice_l166_88;
  reg        [6:0]    _zz_when_ArraySlice_l173_88;
  wire       [5:0]    _zz_when_ArraySlice_l112_88;
  wire                when_ArraySlice_l112_88;
  wire                when_ArraySlice_l113_88;
  wire                when_ArraySlice_l118_88;
  wire                when_ArraySlice_l173_88;
  wire                when_ArraySlice_l165_89;
  wire                when_ArraySlice_l166_89;
  reg        [6:0]    _zz_when_ArraySlice_l173_89;
  wire       [5:0]    _zz_when_ArraySlice_l112_89;
  wire                when_ArraySlice_l112_89;
  wire                when_ArraySlice_l113_89;
  wire                when_ArraySlice_l118_89;
  wire                when_ArraySlice_l173_89;
  wire                when_ArraySlice_l165_90;
  wire                when_ArraySlice_l166_90;
  reg        [6:0]    _zz_when_ArraySlice_l173_90;
  wire       [5:0]    _zz_when_ArraySlice_l112_90;
  wire                when_ArraySlice_l112_90;
  wire                when_ArraySlice_l113_90;
  wire                when_ArraySlice_l118_90;
  wire                when_ArraySlice_l173_90;
  wire                when_ArraySlice_l165_91;
  wire                when_ArraySlice_l166_91;
  reg        [6:0]    _zz_when_ArraySlice_l173_91;
  wire       [5:0]    _zz_when_ArraySlice_l112_91;
  wire                when_ArraySlice_l112_91;
  wire                when_ArraySlice_l113_91;
  wire                when_ArraySlice_l118_91;
  wire                when_ArraySlice_l173_91;
  wire                when_ArraySlice_l165_92;
  wire                when_ArraySlice_l166_92;
  reg        [6:0]    _zz_when_ArraySlice_l173_92;
  wire       [5:0]    _zz_when_ArraySlice_l112_92;
  wire                when_ArraySlice_l112_92;
  wire                when_ArraySlice_l113_92;
  wire                when_ArraySlice_l118_92;
  wire                when_ArraySlice_l173_92;
  wire                when_ArraySlice_l165_93;
  wire                when_ArraySlice_l166_93;
  reg        [6:0]    _zz_when_ArraySlice_l173_93;
  wire       [5:0]    _zz_when_ArraySlice_l112_93;
  wire                when_ArraySlice_l112_93;
  wire                when_ArraySlice_l113_93;
  wire                when_ArraySlice_l118_93;
  wire                when_ArraySlice_l173_93;
  wire                when_ArraySlice_l165_94;
  wire                when_ArraySlice_l166_94;
  reg        [6:0]    _zz_when_ArraySlice_l173_94;
  wire       [5:0]    _zz_when_ArraySlice_l112_94;
  wire                when_ArraySlice_l112_94;
  wire                when_ArraySlice_l113_94;
  wire                when_ArraySlice_l118_94;
  wire                when_ArraySlice_l173_94;
  wire                when_ArraySlice_l165_95;
  wire                when_ArraySlice_l166_95;
  reg        [6:0]    _zz_when_ArraySlice_l173_95;
  wire       [5:0]    _zz_when_ArraySlice_l112_95;
  wire                when_ArraySlice_l112_95;
  wire                when_ArraySlice_l113_95;
  wire                when_ArraySlice_l118_95;
  wire                when_ArraySlice_l173_95;
  wire                when_ArraySlice_l418_3;
  wire                when_ArraySlice_l421_3;
  wire                outputStreamArrayData_3_fire_3;
  wire                when_ArraySlice_l425_3;
  wire                outputStreamArrayData_3_fire_4;
  wire                when_ArraySlice_l436_3;
  reg        [6:0]    _zz_when_ArraySlice_l437_3;
  wire       [5:0]    _zz_when_ArraySlice_l94_11;
  wire                when_ArraySlice_l94_11;
  wire                when_ArraySlice_l95_11;
  wire                when_ArraySlice_l99_11;
  wire                when_ArraySlice_l437_3;
  reg                 debug_0_12 /* verilator public */ ;
  reg                 debug_1_12 /* verilator public */ ;
  reg                 debug_2_12 /* verilator public */ ;
  reg                 debug_3_12 /* verilator public */ ;
  reg                 debug_4_12 /* verilator public */ ;
  reg                 debug_5_12 /* verilator public */ ;
  reg                 debug_6_12 /* verilator public */ ;
  reg                 debug_7_12 /* verilator public */ ;
  wire                when_ArraySlice_l165_96;
  wire                when_ArraySlice_l166_96;
  reg        [6:0]    _zz_when_ArraySlice_l173_96;
  wire       [5:0]    _zz_when_ArraySlice_l112_96;
  wire                when_ArraySlice_l112_96;
  wire                when_ArraySlice_l113_96;
  wire                when_ArraySlice_l118_96;
  wire                when_ArraySlice_l173_96;
  wire                when_ArraySlice_l165_97;
  wire                when_ArraySlice_l166_97;
  reg        [6:0]    _zz_when_ArraySlice_l173_97;
  wire       [5:0]    _zz_when_ArraySlice_l112_97;
  wire                when_ArraySlice_l112_97;
  wire                when_ArraySlice_l113_97;
  wire                when_ArraySlice_l118_97;
  wire                when_ArraySlice_l173_97;
  wire                when_ArraySlice_l165_98;
  wire                when_ArraySlice_l166_98;
  reg        [6:0]    _zz_when_ArraySlice_l173_98;
  wire       [5:0]    _zz_when_ArraySlice_l112_98;
  wire                when_ArraySlice_l112_98;
  wire                when_ArraySlice_l113_98;
  wire                when_ArraySlice_l118_98;
  wire                when_ArraySlice_l173_98;
  wire                when_ArraySlice_l165_99;
  wire                when_ArraySlice_l166_99;
  reg        [6:0]    _zz_when_ArraySlice_l173_99;
  wire       [5:0]    _zz_when_ArraySlice_l112_99;
  wire                when_ArraySlice_l112_99;
  wire                when_ArraySlice_l113_99;
  wire                when_ArraySlice_l118_99;
  wire                when_ArraySlice_l173_99;
  wire                when_ArraySlice_l165_100;
  wire                when_ArraySlice_l166_100;
  reg        [6:0]    _zz_when_ArraySlice_l173_100;
  wire       [5:0]    _zz_when_ArraySlice_l112_100;
  wire                when_ArraySlice_l112_100;
  wire                when_ArraySlice_l113_100;
  wire                when_ArraySlice_l118_100;
  wire                when_ArraySlice_l173_100;
  wire                when_ArraySlice_l165_101;
  wire                when_ArraySlice_l166_101;
  reg        [6:0]    _zz_when_ArraySlice_l173_101;
  wire       [5:0]    _zz_when_ArraySlice_l112_101;
  wire                when_ArraySlice_l112_101;
  wire                when_ArraySlice_l113_101;
  wire                when_ArraySlice_l118_101;
  wire                when_ArraySlice_l173_101;
  wire                when_ArraySlice_l165_102;
  wire                when_ArraySlice_l166_102;
  reg        [6:0]    _zz_when_ArraySlice_l173_102;
  wire       [5:0]    _zz_when_ArraySlice_l112_102;
  wire                when_ArraySlice_l112_102;
  wire                when_ArraySlice_l113_102;
  wire                when_ArraySlice_l118_102;
  wire                when_ArraySlice_l173_102;
  wire                when_ArraySlice_l165_103;
  wire                when_ArraySlice_l166_103;
  reg        [6:0]    _zz_when_ArraySlice_l173_103;
  wire       [5:0]    _zz_when_ArraySlice_l112_103;
  wire                when_ArraySlice_l112_103;
  wire                when_ArraySlice_l113_103;
  wire                when_ArraySlice_l118_103;
  wire                when_ArraySlice_l173_103;
  wire                when_ArraySlice_l444_3;
  wire                outputStreamArrayData_3_fire_5;
  wire                when_ArraySlice_l448_3;
  wire                when_ArraySlice_l434_3;
  wire                outputStreamArrayData_3_fire_6;
  wire                when_ArraySlice_l455_3;
  wire                when_ArraySlice_l373_4;
  wire                when_ArraySlice_l374_4;
  wire       [5:0]    _zz_outputStreamArrayData_4_valid;
  wire                _zz_io_pop_ready_4;
  wire       [63:0]   _zz_7;
  wire                when_ArraySlice_l379_4;
  wire                outputStreamArrayData_4_fire;
  wire                when_ArraySlice_l380_4;
  wire                when_ArraySlice_l381_4;
  wire                when_ArraySlice_l384_4;
  wire                outputStreamArrayData_4_fire_1;
  wire                when_ArraySlice_l389_4;
  wire                when_ArraySlice_l390_4;
  reg        [6:0]    _zz_when_ArraySlice_l392_4;
  wire       [5:0]    _zz_when_ArraySlice_l94_12;
  wire                when_ArraySlice_l94_12;
  wire                when_ArraySlice_l95_12;
  wire                when_ArraySlice_l99_12;
  wire                when_ArraySlice_l392_4;
  reg                 debug_0_13 /* verilator public */ ;
  reg                 debug_1_13 /* verilator public */ ;
  reg                 debug_2_13 /* verilator public */ ;
  reg                 debug_3_13 /* verilator public */ ;
  reg                 debug_4_13 /* verilator public */ ;
  reg                 debug_5_13 /* verilator public */ ;
  reg                 debug_6_13 /* verilator public */ ;
  reg                 debug_7_13 /* verilator public */ ;
  wire                when_ArraySlice_l165_104;
  wire                when_ArraySlice_l166_104;
  reg        [6:0]    _zz_when_ArraySlice_l173_104;
  wire       [5:0]    _zz_when_ArraySlice_l112_104;
  wire                when_ArraySlice_l112_104;
  wire                when_ArraySlice_l113_104;
  wire                when_ArraySlice_l118_104;
  wire                when_ArraySlice_l173_104;
  wire                when_ArraySlice_l165_105;
  wire                when_ArraySlice_l166_105;
  reg        [6:0]    _zz_when_ArraySlice_l173_105;
  wire       [5:0]    _zz_when_ArraySlice_l112_105;
  wire                when_ArraySlice_l112_105;
  wire                when_ArraySlice_l113_105;
  wire                when_ArraySlice_l118_105;
  wire                when_ArraySlice_l173_105;
  wire                when_ArraySlice_l165_106;
  wire                when_ArraySlice_l166_106;
  reg        [6:0]    _zz_when_ArraySlice_l173_106;
  wire       [5:0]    _zz_when_ArraySlice_l112_106;
  wire                when_ArraySlice_l112_106;
  wire                when_ArraySlice_l113_106;
  wire                when_ArraySlice_l118_106;
  wire                when_ArraySlice_l173_106;
  wire                when_ArraySlice_l165_107;
  wire                when_ArraySlice_l166_107;
  reg        [6:0]    _zz_when_ArraySlice_l173_107;
  wire       [5:0]    _zz_when_ArraySlice_l112_107;
  wire                when_ArraySlice_l112_107;
  wire                when_ArraySlice_l113_107;
  wire                when_ArraySlice_l118_107;
  wire                when_ArraySlice_l173_107;
  wire                when_ArraySlice_l165_108;
  wire                when_ArraySlice_l166_108;
  reg        [6:0]    _zz_when_ArraySlice_l173_108;
  wire       [5:0]    _zz_when_ArraySlice_l112_108;
  wire                when_ArraySlice_l112_108;
  wire                when_ArraySlice_l113_108;
  wire                when_ArraySlice_l118_108;
  wire                when_ArraySlice_l173_108;
  wire                when_ArraySlice_l165_109;
  wire                when_ArraySlice_l166_109;
  reg        [6:0]    _zz_when_ArraySlice_l173_109;
  wire       [5:0]    _zz_when_ArraySlice_l112_109;
  wire                when_ArraySlice_l112_109;
  wire                when_ArraySlice_l113_109;
  wire                when_ArraySlice_l118_109;
  wire                when_ArraySlice_l173_109;
  wire                when_ArraySlice_l165_110;
  wire                when_ArraySlice_l166_110;
  reg        [6:0]    _zz_when_ArraySlice_l173_110;
  wire       [5:0]    _zz_when_ArraySlice_l112_110;
  wire                when_ArraySlice_l112_110;
  wire                when_ArraySlice_l113_110;
  wire                when_ArraySlice_l118_110;
  wire                when_ArraySlice_l173_110;
  wire                when_ArraySlice_l165_111;
  wire                when_ArraySlice_l166_111;
  reg        [6:0]    _zz_when_ArraySlice_l173_111;
  wire       [5:0]    _zz_when_ArraySlice_l112_111;
  wire                when_ArraySlice_l112_111;
  wire                when_ArraySlice_l113_111;
  wire                when_ArraySlice_l118_111;
  wire                when_ArraySlice_l173_111;
  wire                when_ArraySlice_l398_4;
  wire                when_ArraySlice_l401_4;
  wire                when_ArraySlice_l405_4;
  wire                when_ArraySlice_l409_4;
  wire                outputStreamArrayData_4_fire_2;
  wire                when_ArraySlice_l410_4;
  reg        [6:0]    _zz_when_ArraySlice_l412_4;
  wire       [5:0]    _zz_when_ArraySlice_l94_13;
  wire                when_ArraySlice_l94_13;
  wire                when_ArraySlice_l95_13;
  wire                when_ArraySlice_l99_13;
  wire                when_ArraySlice_l412_4;
  reg                 debug_0_14 /* verilator public */ ;
  reg                 debug_1_14 /* verilator public */ ;
  reg                 debug_2_14 /* verilator public */ ;
  reg                 debug_3_14 /* verilator public */ ;
  reg                 debug_4_14 /* verilator public */ ;
  reg                 debug_5_14 /* verilator public */ ;
  reg                 debug_6_14 /* verilator public */ ;
  reg                 debug_7_14 /* verilator public */ ;
  wire                when_ArraySlice_l165_112;
  wire                when_ArraySlice_l166_112;
  reg        [6:0]    _zz_when_ArraySlice_l173_112;
  wire       [5:0]    _zz_when_ArraySlice_l112_112;
  wire                when_ArraySlice_l112_112;
  wire                when_ArraySlice_l113_112;
  wire                when_ArraySlice_l118_112;
  wire                when_ArraySlice_l173_112;
  wire                when_ArraySlice_l165_113;
  wire                when_ArraySlice_l166_113;
  reg        [6:0]    _zz_when_ArraySlice_l173_113;
  wire       [5:0]    _zz_when_ArraySlice_l112_113;
  wire                when_ArraySlice_l112_113;
  wire                when_ArraySlice_l113_113;
  wire                when_ArraySlice_l118_113;
  wire                when_ArraySlice_l173_113;
  wire                when_ArraySlice_l165_114;
  wire                when_ArraySlice_l166_114;
  reg        [6:0]    _zz_when_ArraySlice_l173_114;
  wire       [5:0]    _zz_when_ArraySlice_l112_114;
  wire                when_ArraySlice_l112_114;
  wire                when_ArraySlice_l113_114;
  wire                when_ArraySlice_l118_114;
  wire                when_ArraySlice_l173_114;
  wire                when_ArraySlice_l165_115;
  wire                when_ArraySlice_l166_115;
  reg        [6:0]    _zz_when_ArraySlice_l173_115;
  wire       [5:0]    _zz_when_ArraySlice_l112_115;
  wire                when_ArraySlice_l112_115;
  wire                when_ArraySlice_l113_115;
  wire                when_ArraySlice_l118_115;
  wire                when_ArraySlice_l173_115;
  wire                when_ArraySlice_l165_116;
  wire                when_ArraySlice_l166_116;
  reg        [6:0]    _zz_when_ArraySlice_l173_116;
  wire       [5:0]    _zz_when_ArraySlice_l112_116;
  wire                when_ArraySlice_l112_116;
  wire                when_ArraySlice_l113_116;
  wire                when_ArraySlice_l118_116;
  wire                when_ArraySlice_l173_116;
  wire                when_ArraySlice_l165_117;
  wire                when_ArraySlice_l166_117;
  reg        [6:0]    _zz_when_ArraySlice_l173_117;
  wire       [5:0]    _zz_when_ArraySlice_l112_117;
  wire                when_ArraySlice_l112_117;
  wire                when_ArraySlice_l113_117;
  wire                when_ArraySlice_l118_117;
  wire                when_ArraySlice_l173_117;
  wire                when_ArraySlice_l165_118;
  wire                when_ArraySlice_l166_118;
  reg        [6:0]    _zz_when_ArraySlice_l173_118;
  wire       [5:0]    _zz_when_ArraySlice_l112_118;
  wire                when_ArraySlice_l112_118;
  wire                when_ArraySlice_l113_118;
  wire                when_ArraySlice_l118_118;
  wire                when_ArraySlice_l173_118;
  wire                when_ArraySlice_l165_119;
  wire                when_ArraySlice_l166_119;
  reg        [6:0]    _zz_when_ArraySlice_l173_119;
  wire       [5:0]    _zz_when_ArraySlice_l112_119;
  wire                when_ArraySlice_l112_119;
  wire                when_ArraySlice_l113_119;
  wire                when_ArraySlice_l118_119;
  wire                when_ArraySlice_l173_119;
  wire                when_ArraySlice_l418_4;
  wire                when_ArraySlice_l421_4;
  wire                outputStreamArrayData_4_fire_3;
  wire                when_ArraySlice_l425_4;
  wire                outputStreamArrayData_4_fire_4;
  wire                when_ArraySlice_l436_4;
  reg        [6:0]    _zz_when_ArraySlice_l437_4;
  wire       [5:0]    _zz_when_ArraySlice_l94_14;
  wire                when_ArraySlice_l94_14;
  wire                when_ArraySlice_l95_14;
  wire                when_ArraySlice_l99_14;
  wire                when_ArraySlice_l437_4;
  reg                 debug_0_15 /* verilator public */ ;
  reg                 debug_1_15 /* verilator public */ ;
  reg                 debug_2_15 /* verilator public */ ;
  reg                 debug_3_15 /* verilator public */ ;
  reg                 debug_4_15 /* verilator public */ ;
  reg                 debug_5_15 /* verilator public */ ;
  reg                 debug_6_15 /* verilator public */ ;
  reg                 debug_7_15 /* verilator public */ ;
  wire                when_ArraySlice_l165_120;
  wire                when_ArraySlice_l166_120;
  reg        [6:0]    _zz_when_ArraySlice_l173_120;
  wire       [5:0]    _zz_when_ArraySlice_l112_120;
  wire                when_ArraySlice_l112_120;
  wire                when_ArraySlice_l113_120;
  wire                when_ArraySlice_l118_120;
  wire                when_ArraySlice_l173_120;
  wire                when_ArraySlice_l165_121;
  wire                when_ArraySlice_l166_121;
  reg        [6:0]    _zz_when_ArraySlice_l173_121;
  wire       [5:0]    _zz_when_ArraySlice_l112_121;
  wire                when_ArraySlice_l112_121;
  wire                when_ArraySlice_l113_121;
  wire                when_ArraySlice_l118_121;
  wire                when_ArraySlice_l173_121;
  wire                when_ArraySlice_l165_122;
  wire                when_ArraySlice_l166_122;
  reg        [6:0]    _zz_when_ArraySlice_l173_122;
  wire       [5:0]    _zz_when_ArraySlice_l112_122;
  wire                when_ArraySlice_l112_122;
  wire                when_ArraySlice_l113_122;
  wire                when_ArraySlice_l118_122;
  wire                when_ArraySlice_l173_122;
  wire                when_ArraySlice_l165_123;
  wire                when_ArraySlice_l166_123;
  reg        [6:0]    _zz_when_ArraySlice_l173_123;
  wire       [5:0]    _zz_when_ArraySlice_l112_123;
  wire                when_ArraySlice_l112_123;
  wire                when_ArraySlice_l113_123;
  wire                when_ArraySlice_l118_123;
  wire                when_ArraySlice_l173_123;
  wire                when_ArraySlice_l165_124;
  wire                when_ArraySlice_l166_124;
  reg        [6:0]    _zz_when_ArraySlice_l173_124;
  wire       [5:0]    _zz_when_ArraySlice_l112_124;
  wire                when_ArraySlice_l112_124;
  wire                when_ArraySlice_l113_124;
  wire                when_ArraySlice_l118_124;
  wire                when_ArraySlice_l173_124;
  wire                when_ArraySlice_l165_125;
  wire                when_ArraySlice_l166_125;
  reg        [6:0]    _zz_when_ArraySlice_l173_125;
  wire       [5:0]    _zz_when_ArraySlice_l112_125;
  wire                when_ArraySlice_l112_125;
  wire                when_ArraySlice_l113_125;
  wire                when_ArraySlice_l118_125;
  wire                when_ArraySlice_l173_125;
  wire                when_ArraySlice_l165_126;
  wire                when_ArraySlice_l166_126;
  reg        [6:0]    _zz_when_ArraySlice_l173_126;
  wire       [5:0]    _zz_when_ArraySlice_l112_126;
  wire                when_ArraySlice_l112_126;
  wire                when_ArraySlice_l113_126;
  wire                when_ArraySlice_l118_126;
  wire                when_ArraySlice_l173_126;
  wire                when_ArraySlice_l165_127;
  wire                when_ArraySlice_l166_127;
  reg        [6:0]    _zz_when_ArraySlice_l173_127;
  wire       [5:0]    _zz_when_ArraySlice_l112_127;
  wire                when_ArraySlice_l112_127;
  wire                when_ArraySlice_l113_127;
  wire                when_ArraySlice_l118_127;
  wire                when_ArraySlice_l173_127;
  wire                when_ArraySlice_l444_4;
  wire                outputStreamArrayData_4_fire_5;
  wire                when_ArraySlice_l448_4;
  wire                when_ArraySlice_l434_4;
  wire                outputStreamArrayData_4_fire_6;
  wire                when_ArraySlice_l455_4;
  wire                when_ArraySlice_l373_5;
  wire                when_ArraySlice_l374_5;
  wire       [5:0]    _zz_outputStreamArrayData_5_valid;
  wire                _zz_io_pop_ready_5;
  wire       [63:0]   _zz_8;
  wire                when_ArraySlice_l379_5;
  wire                outputStreamArrayData_5_fire;
  wire                when_ArraySlice_l380_5;
  wire                when_ArraySlice_l381_5;
  wire                when_ArraySlice_l384_5;
  wire                outputStreamArrayData_5_fire_1;
  wire                when_ArraySlice_l389_5;
  wire                when_ArraySlice_l390_5;
  reg        [6:0]    _zz_when_ArraySlice_l392_5;
  wire       [5:0]    _zz_when_ArraySlice_l94_15;
  wire                when_ArraySlice_l94_15;
  wire                when_ArraySlice_l95_15;
  wire                when_ArraySlice_l99_15;
  wire                when_ArraySlice_l392_5;
  reg                 debug_0_16 /* verilator public */ ;
  reg                 debug_1_16 /* verilator public */ ;
  reg                 debug_2_16 /* verilator public */ ;
  reg                 debug_3_16 /* verilator public */ ;
  reg                 debug_4_16 /* verilator public */ ;
  reg                 debug_5_16 /* verilator public */ ;
  reg                 debug_6_16 /* verilator public */ ;
  reg                 debug_7_16 /* verilator public */ ;
  wire                when_ArraySlice_l165_128;
  wire                when_ArraySlice_l166_128;
  reg        [6:0]    _zz_when_ArraySlice_l173_128;
  wire       [5:0]    _zz_when_ArraySlice_l112_128;
  wire                when_ArraySlice_l112_128;
  wire                when_ArraySlice_l113_128;
  wire                when_ArraySlice_l118_128;
  wire                when_ArraySlice_l173_128;
  wire                when_ArraySlice_l165_129;
  wire                when_ArraySlice_l166_129;
  reg        [6:0]    _zz_when_ArraySlice_l173_129;
  wire       [5:0]    _zz_when_ArraySlice_l112_129;
  wire                when_ArraySlice_l112_129;
  wire                when_ArraySlice_l113_129;
  wire                when_ArraySlice_l118_129;
  wire                when_ArraySlice_l173_129;
  wire                when_ArraySlice_l165_130;
  wire                when_ArraySlice_l166_130;
  reg        [6:0]    _zz_when_ArraySlice_l173_130;
  wire       [5:0]    _zz_when_ArraySlice_l112_130;
  wire                when_ArraySlice_l112_130;
  wire                when_ArraySlice_l113_130;
  wire                when_ArraySlice_l118_130;
  wire                when_ArraySlice_l173_130;
  wire                when_ArraySlice_l165_131;
  wire                when_ArraySlice_l166_131;
  reg        [6:0]    _zz_when_ArraySlice_l173_131;
  wire       [5:0]    _zz_when_ArraySlice_l112_131;
  wire                when_ArraySlice_l112_131;
  wire                when_ArraySlice_l113_131;
  wire                when_ArraySlice_l118_131;
  wire                when_ArraySlice_l173_131;
  wire                when_ArraySlice_l165_132;
  wire                when_ArraySlice_l166_132;
  reg        [6:0]    _zz_when_ArraySlice_l173_132;
  wire       [5:0]    _zz_when_ArraySlice_l112_132;
  wire                when_ArraySlice_l112_132;
  wire                when_ArraySlice_l113_132;
  wire                when_ArraySlice_l118_132;
  wire                when_ArraySlice_l173_132;
  wire                when_ArraySlice_l165_133;
  wire                when_ArraySlice_l166_133;
  reg        [6:0]    _zz_when_ArraySlice_l173_133;
  wire       [5:0]    _zz_when_ArraySlice_l112_133;
  wire                when_ArraySlice_l112_133;
  wire                when_ArraySlice_l113_133;
  wire                when_ArraySlice_l118_133;
  wire                when_ArraySlice_l173_133;
  wire                when_ArraySlice_l165_134;
  wire                when_ArraySlice_l166_134;
  reg        [6:0]    _zz_when_ArraySlice_l173_134;
  wire       [5:0]    _zz_when_ArraySlice_l112_134;
  wire                when_ArraySlice_l112_134;
  wire                when_ArraySlice_l113_134;
  wire                when_ArraySlice_l118_134;
  wire                when_ArraySlice_l173_134;
  wire                when_ArraySlice_l165_135;
  wire                when_ArraySlice_l166_135;
  reg        [6:0]    _zz_when_ArraySlice_l173_135;
  wire       [5:0]    _zz_when_ArraySlice_l112_135;
  wire                when_ArraySlice_l112_135;
  wire                when_ArraySlice_l113_135;
  wire                when_ArraySlice_l118_135;
  wire                when_ArraySlice_l173_135;
  wire                when_ArraySlice_l398_5;
  wire                when_ArraySlice_l401_5;
  wire                when_ArraySlice_l405_5;
  wire                when_ArraySlice_l409_5;
  wire                outputStreamArrayData_5_fire_2;
  wire                when_ArraySlice_l410_5;
  reg        [6:0]    _zz_when_ArraySlice_l412_5;
  wire       [5:0]    _zz_when_ArraySlice_l94_16;
  wire                when_ArraySlice_l94_16;
  wire                when_ArraySlice_l95_16;
  wire                when_ArraySlice_l99_16;
  wire                when_ArraySlice_l412_5;
  reg                 debug_0_17 /* verilator public */ ;
  reg                 debug_1_17 /* verilator public */ ;
  reg                 debug_2_17 /* verilator public */ ;
  reg                 debug_3_17 /* verilator public */ ;
  reg                 debug_4_17 /* verilator public */ ;
  reg                 debug_5_17 /* verilator public */ ;
  reg                 debug_6_17 /* verilator public */ ;
  reg                 debug_7_17 /* verilator public */ ;
  wire                when_ArraySlice_l165_136;
  wire                when_ArraySlice_l166_136;
  reg        [6:0]    _zz_when_ArraySlice_l173_136;
  wire       [5:0]    _zz_when_ArraySlice_l112_136;
  wire                when_ArraySlice_l112_136;
  wire                when_ArraySlice_l113_136;
  wire                when_ArraySlice_l118_136;
  wire                when_ArraySlice_l173_136;
  wire                when_ArraySlice_l165_137;
  wire                when_ArraySlice_l166_137;
  reg        [6:0]    _zz_when_ArraySlice_l173_137;
  wire       [5:0]    _zz_when_ArraySlice_l112_137;
  wire                when_ArraySlice_l112_137;
  wire                when_ArraySlice_l113_137;
  wire                when_ArraySlice_l118_137;
  wire                when_ArraySlice_l173_137;
  wire                when_ArraySlice_l165_138;
  wire                when_ArraySlice_l166_138;
  reg        [6:0]    _zz_when_ArraySlice_l173_138;
  wire       [5:0]    _zz_when_ArraySlice_l112_138;
  wire                when_ArraySlice_l112_138;
  wire                when_ArraySlice_l113_138;
  wire                when_ArraySlice_l118_138;
  wire                when_ArraySlice_l173_138;
  wire                when_ArraySlice_l165_139;
  wire                when_ArraySlice_l166_139;
  reg        [6:0]    _zz_when_ArraySlice_l173_139;
  wire       [5:0]    _zz_when_ArraySlice_l112_139;
  wire                when_ArraySlice_l112_139;
  wire                when_ArraySlice_l113_139;
  wire                when_ArraySlice_l118_139;
  wire                when_ArraySlice_l173_139;
  wire                when_ArraySlice_l165_140;
  wire                when_ArraySlice_l166_140;
  reg        [6:0]    _zz_when_ArraySlice_l173_140;
  wire       [5:0]    _zz_when_ArraySlice_l112_140;
  wire                when_ArraySlice_l112_140;
  wire                when_ArraySlice_l113_140;
  wire                when_ArraySlice_l118_140;
  wire                when_ArraySlice_l173_140;
  wire                when_ArraySlice_l165_141;
  wire                when_ArraySlice_l166_141;
  reg        [6:0]    _zz_when_ArraySlice_l173_141;
  wire       [5:0]    _zz_when_ArraySlice_l112_141;
  wire                when_ArraySlice_l112_141;
  wire                when_ArraySlice_l113_141;
  wire                when_ArraySlice_l118_141;
  wire                when_ArraySlice_l173_141;
  wire                when_ArraySlice_l165_142;
  wire                when_ArraySlice_l166_142;
  reg        [6:0]    _zz_when_ArraySlice_l173_142;
  wire       [5:0]    _zz_when_ArraySlice_l112_142;
  wire                when_ArraySlice_l112_142;
  wire                when_ArraySlice_l113_142;
  wire                when_ArraySlice_l118_142;
  wire                when_ArraySlice_l173_142;
  wire                when_ArraySlice_l165_143;
  wire                when_ArraySlice_l166_143;
  reg        [6:0]    _zz_when_ArraySlice_l173_143;
  wire       [5:0]    _zz_when_ArraySlice_l112_143;
  wire                when_ArraySlice_l112_143;
  wire                when_ArraySlice_l113_143;
  wire                when_ArraySlice_l118_143;
  wire                when_ArraySlice_l173_143;
  wire                when_ArraySlice_l418_5;
  wire                when_ArraySlice_l421_5;
  wire                outputStreamArrayData_5_fire_3;
  wire                when_ArraySlice_l425_5;
  wire                outputStreamArrayData_5_fire_4;
  wire                when_ArraySlice_l436_5;
  reg        [6:0]    _zz_when_ArraySlice_l437_5;
  wire       [5:0]    _zz_when_ArraySlice_l94_17;
  wire                when_ArraySlice_l94_17;
  wire                when_ArraySlice_l95_17;
  wire                when_ArraySlice_l99_17;
  wire                when_ArraySlice_l437_5;
  reg                 debug_0_18 /* verilator public */ ;
  reg                 debug_1_18 /* verilator public */ ;
  reg                 debug_2_18 /* verilator public */ ;
  reg                 debug_3_18 /* verilator public */ ;
  reg                 debug_4_18 /* verilator public */ ;
  reg                 debug_5_18 /* verilator public */ ;
  reg                 debug_6_18 /* verilator public */ ;
  reg                 debug_7_18 /* verilator public */ ;
  wire                when_ArraySlice_l165_144;
  wire                when_ArraySlice_l166_144;
  reg        [6:0]    _zz_when_ArraySlice_l173_144;
  wire       [5:0]    _zz_when_ArraySlice_l112_144;
  wire                when_ArraySlice_l112_144;
  wire                when_ArraySlice_l113_144;
  wire                when_ArraySlice_l118_144;
  wire                when_ArraySlice_l173_144;
  wire                when_ArraySlice_l165_145;
  wire                when_ArraySlice_l166_145;
  reg        [6:0]    _zz_when_ArraySlice_l173_145;
  wire       [5:0]    _zz_when_ArraySlice_l112_145;
  wire                when_ArraySlice_l112_145;
  wire                when_ArraySlice_l113_145;
  wire                when_ArraySlice_l118_145;
  wire                when_ArraySlice_l173_145;
  wire                when_ArraySlice_l165_146;
  wire                when_ArraySlice_l166_146;
  reg        [6:0]    _zz_when_ArraySlice_l173_146;
  wire       [5:0]    _zz_when_ArraySlice_l112_146;
  wire                when_ArraySlice_l112_146;
  wire                when_ArraySlice_l113_146;
  wire                when_ArraySlice_l118_146;
  wire                when_ArraySlice_l173_146;
  wire                when_ArraySlice_l165_147;
  wire                when_ArraySlice_l166_147;
  reg        [6:0]    _zz_when_ArraySlice_l173_147;
  wire       [5:0]    _zz_when_ArraySlice_l112_147;
  wire                when_ArraySlice_l112_147;
  wire                when_ArraySlice_l113_147;
  wire                when_ArraySlice_l118_147;
  wire                when_ArraySlice_l173_147;
  wire                when_ArraySlice_l165_148;
  wire                when_ArraySlice_l166_148;
  reg        [6:0]    _zz_when_ArraySlice_l173_148;
  wire       [5:0]    _zz_when_ArraySlice_l112_148;
  wire                when_ArraySlice_l112_148;
  wire                when_ArraySlice_l113_148;
  wire                when_ArraySlice_l118_148;
  wire                when_ArraySlice_l173_148;
  wire                when_ArraySlice_l165_149;
  wire                when_ArraySlice_l166_149;
  reg        [6:0]    _zz_when_ArraySlice_l173_149;
  wire       [5:0]    _zz_when_ArraySlice_l112_149;
  wire                when_ArraySlice_l112_149;
  wire                when_ArraySlice_l113_149;
  wire                when_ArraySlice_l118_149;
  wire                when_ArraySlice_l173_149;
  wire                when_ArraySlice_l165_150;
  wire                when_ArraySlice_l166_150;
  reg        [6:0]    _zz_when_ArraySlice_l173_150;
  wire       [5:0]    _zz_when_ArraySlice_l112_150;
  wire                when_ArraySlice_l112_150;
  wire                when_ArraySlice_l113_150;
  wire                when_ArraySlice_l118_150;
  wire                when_ArraySlice_l173_150;
  wire                when_ArraySlice_l165_151;
  wire                when_ArraySlice_l166_151;
  reg        [6:0]    _zz_when_ArraySlice_l173_151;
  wire       [5:0]    _zz_when_ArraySlice_l112_151;
  wire                when_ArraySlice_l112_151;
  wire                when_ArraySlice_l113_151;
  wire                when_ArraySlice_l118_151;
  wire                when_ArraySlice_l173_151;
  wire                when_ArraySlice_l444_5;
  wire                outputStreamArrayData_5_fire_5;
  wire                when_ArraySlice_l448_5;
  wire                when_ArraySlice_l434_5;
  wire                outputStreamArrayData_5_fire_6;
  wire                when_ArraySlice_l455_5;
  wire                when_ArraySlice_l373_6;
  wire                when_ArraySlice_l374_6;
  wire       [5:0]    _zz_outputStreamArrayData_6_valid;
  wire                _zz_io_pop_ready_6;
  wire       [63:0]   _zz_9;
  wire                when_ArraySlice_l379_6;
  wire                outputStreamArrayData_6_fire;
  wire                when_ArraySlice_l380_6;
  wire                when_ArraySlice_l381_6;
  wire                when_ArraySlice_l384_6;
  wire                outputStreamArrayData_6_fire_1;
  wire                when_ArraySlice_l389_6;
  wire                when_ArraySlice_l390_6;
  reg        [6:0]    _zz_when_ArraySlice_l392_6;
  wire       [5:0]    _zz_when_ArraySlice_l94_18;
  wire                when_ArraySlice_l94_18;
  wire                when_ArraySlice_l95_18;
  wire                when_ArraySlice_l99_18;
  wire                when_ArraySlice_l392_6;
  reg                 debug_0_19 /* verilator public */ ;
  reg                 debug_1_19 /* verilator public */ ;
  reg                 debug_2_19 /* verilator public */ ;
  reg                 debug_3_19 /* verilator public */ ;
  reg                 debug_4_19 /* verilator public */ ;
  reg                 debug_5_19 /* verilator public */ ;
  reg                 debug_6_19 /* verilator public */ ;
  reg                 debug_7_19 /* verilator public */ ;
  wire                when_ArraySlice_l165_152;
  wire                when_ArraySlice_l166_152;
  reg        [6:0]    _zz_when_ArraySlice_l173_152;
  wire       [5:0]    _zz_when_ArraySlice_l112_152;
  wire                when_ArraySlice_l112_152;
  wire                when_ArraySlice_l113_152;
  wire                when_ArraySlice_l118_152;
  wire                when_ArraySlice_l173_152;
  wire                when_ArraySlice_l165_153;
  wire                when_ArraySlice_l166_153;
  reg        [6:0]    _zz_when_ArraySlice_l173_153;
  wire       [5:0]    _zz_when_ArraySlice_l112_153;
  wire                when_ArraySlice_l112_153;
  wire                when_ArraySlice_l113_153;
  wire                when_ArraySlice_l118_153;
  wire                when_ArraySlice_l173_153;
  wire                when_ArraySlice_l165_154;
  wire                when_ArraySlice_l166_154;
  reg        [6:0]    _zz_when_ArraySlice_l173_154;
  wire       [5:0]    _zz_when_ArraySlice_l112_154;
  wire                when_ArraySlice_l112_154;
  wire                when_ArraySlice_l113_154;
  wire                when_ArraySlice_l118_154;
  wire                when_ArraySlice_l173_154;
  wire                when_ArraySlice_l165_155;
  wire                when_ArraySlice_l166_155;
  reg        [6:0]    _zz_when_ArraySlice_l173_155;
  wire       [5:0]    _zz_when_ArraySlice_l112_155;
  wire                when_ArraySlice_l112_155;
  wire                when_ArraySlice_l113_155;
  wire                when_ArraySlice_l118_155;
  wire                when_ArraySlice_l173_155;
  wire                when_ArraySlice_l165_156;
  wire                when_ArraySlice_l166_156;
  reg        [6:0]    _zz_when_ArraySlice_l173_156;
  wire       [5:0]    _zz_when_ArraySlice_l112_156;
  wire                when_ArraySlice_l112_156;
  wire                when_ArraySlice_l113_156;
  wire                when_ArraySlice_l118_156;
  wire                when_ArraySlice_l173_156;
  wire                when_ArraySlice_l165_157;
  wire                when_ArraySlice_l166_157;
  reg        [6:0]    _zz_when_ArraySlice_l173_157;
  wire       [5:0]    _zz_when_ArraySlice_l112_157;
  wire                when_ArraySlice_l112_157;
  wire                when_ArraySlice_l113_157;
  wire                when_ArraySlice_l118_157;
  wire                when_ArraySlice_l173_157;
  wire                when_ArraySlice_l165_158;
  wire                when_ArraySlice_l166_158;
  reg        [6:0]    _zz_when_ArraySlice_l173_158;
  wire       [5:0]    _zz_when_ArraySlice_l112_158;
  wire                when_ArraySlice_l112_158;
  wire                when_ArraySlice_l113_158;
  wire                when_ArraySlice_l118_158;
  wire                when_ArraySlice_l173_158;
  wire                when_ArraySlice_l165_159;
  wire                when_ArraySlice_l166_159;
  reg        [6:0]    _zz_when_ArraySlice_l173_159;
  wire       [5:0]    _zz_when_ArraySlice_l112_159;
  wire                when_ArraySlice_l112_159;
  wire                when_ArraySlice_l113_159;
  wire                when_ArraySlice_l118_159;
  wire                when_ArraySlice_l173_159;
  wire                when_ArraySlice_l398_6;
  wire                when_ArraySlice_l401_6;
  wire                when_ArraySlice_l405_6;
  wire                when_ArraySlice_l409_6;
  wire                outputStreamArrayData_6_fire_2;
  wire                when_ArraySlice_l410_6;
  reg        [6:0]    _zz_when_ArraySlice_l412_6;
  wire       [5:0]    _zz_when_ArraySlice_l94_19;
  wire                when_ArraySlice_l94_19;
  wire                when_ArraySlice_l95_19;
  wire                when_ArraySlice_l99_19;
  wire                when_ArraySlice_l412_6;
  reg                 debug_0_20 /* verilator public */ ;
  reg                 debug_1_20 /* verilator public */ ;
  reg                 debug_2_20 /* verilator public */ ;
  reg                 debug_3_20 /* verilator public */ ;
  reg                 debug_4_20 /* verilator public */ ;
  reg                 debug_5_20 /* verilator public */ ;
  reg                 debug_6_20 /* verilator public */ ;
  reg                 debug_7_20 /* verilator public */ ;
  wire                when_ArraySlice_l165_160;
  wire                when_ArraySlice_l166_160;
  reg        [6:0]    _zz_when_ArraySlice_l173_160;
  wire       [5:0]    _zz_when_ArraySlice_l112_160;
  wire                when_ArraySlice_l112_160;
  wire                when_ArraySlice_l113_160;
  wire                when_ArraySlice_l118_160;
  wire                when_ArraySlice_l173_160;
  wire                when_ArraySlice_l165_161;
  wire                when_ArraySlice_l166_161;
  reg        [6:0]    _zz_when_ArraySlice_l173_161;
  wire       [5:0]    _zz_when_ArraySlice_l112_161;
  wire                when_ArraySlice_l112_161;
  wire                when_ArraySlice_l113_161;
  wire                when_ArraySlice_l118_161;
  wire                when_ArraySlice_l173_161;
  wire                when_ArraySlice_l165_162;
  wire                when_ArraySlice_l166_162;
  reg        [6:0]    _zz_when_ArraySlice_l173_162;
  wire       [5:0]    _zz_when_ArraySlice_l112_162;
  wire                when_ArraySlice_l112_162;
  wire                when_ArraySlice_l113_162;
  wire                when_ArraySlice_l118_162;
  wire                when_ArraySlice_l173_162;
  wire                when_ArraySlice_l165_163;
  wire                when_ArraySlice_l166_163;
  reg        [6:0]    _zz_when_ArraySlice_l173_163;
  wire       [5:0]    _zz_when_ArraySlice_l112_163;
  wire                when_ArraySlice_l112_163;
  wire                when_ArraySlice_l113_163;
  wire                when_ArraySlice_l118_163;
  wire                when_ArraySlice_l173_163;
  wire                when_ArraySlice_l165_164;
  wire                when_ArraySlice_l166_164;
  reg        [6:0]    _zz_when_ArraySlice_l173_164;
  wire       [5:0]    _zz_when_ArraySlice_l112_164;
  wire                when_ArraySlice_l112_164;
  wire                when_ArraySlice_l113_164;
  wire                when_ArraySlice_l118_164;
  wire                when_ArraySlice_l173_164;
  wire                when_ArraySlice_l165_165;
  wire                when_ArraySlice_l166_165;
  reg        [6:0]    _zz_when_ArraySlice_l173_165;
  wire       [5:0]    _zz_when_ArraySlice_l112_165;
  wire                when_ArraySlice_l112_165;
  wire                when_ArraySlice_l113_165;
  wire                when_ArraySlice_l118_165;
  wire                when_ArraySlice_l173_165;
  wire                when_ArraySlice_l165_166;
  wire                when_ArraySlice_l166_166;
  reg        [6:0]    _zz_when_ArraySlice_l173_166;
  wire       [5:0]    _zz_when_ArraySlice_l112_166;
  wire                when_ArraySlice_l112_166;
  wire                when_ArraySlice_l113_166;
  wire                when_ArraySlice_l118_166;
  wire                when_ArraySlice_l173_166;
  wire                when_ArraySlice_l165_167;
  wire                when_ArraySlice_l166_167;
  reg        [6:0]    _zz_when_ArraySlice_l173_167;
  wire       [5:0]    _zz_when_ArraySlice_l112_167;
  wire                when_ArraySlice_l112_167;
  wire                when_ArraySlice_l113_167;
  wire                when_ArraySlice_l118_167;
  wire                when_ArraySlice_l173_167;
  wire                when_ArraySlice_l418_6;
  wire                when_ArraySlice_l421_6;
  wire                outputStreamArrayData_6_fire_3;
  wire                when_ArraySlice_l425_6;
  wire                outputStreamArrayData_6_fire_4;
  wire                when_ArraySlice_l436_6;
  reg        [6:0]    _zz_when_ArraySlice_l437_6;
  wire       [5:0]    _zz_when_ArraySlice_l94_20;
  wire                when_ArraySlice_l94_20;
  wire                when_ArraySlice_l95_20;
  wire                when_ArraySlice_l99_20;
  wire                when_ArraySlice_l437_6;
  reg                 debug_0_21 /* verilator public */ ;
  reg                 debug_1_21 /* verilator public */ ;
  reg                 debug_2_21 /* verilator public */ ;
  reg                 debug_3_21 /* verilator public */ ;
  reg                 debug_4_21 /* verilator public */ ;
  reg                 debug_5_21 /* verilator public */ ;
  reg                 debug_6_21 /* verilator public */ ;
  reg                 debug_7_21 /* verilator public */ ;
  wire                when_ArraySlice_l165_168;
  wire                when_ArraySlice_l166_168;
  reg        [6:0]    _zz_when_ArraySlice_l173_168;
  wire       [5:0]    _zz_when_ArraySlice_l112_168;
  wire                when_ArraySlice_l112_168;
  wire                when_ArraySlice_l113_168;
  wire                when_ArraySlice_l118_168;
  wire                when_ArraySlice_l173_168;
  wire                when_ArraySlice_l165_169;
  wire                when_ArraySlice_l166_169;
  reg        [6:0]    _zz_when_ArraySlice_l173_169;
  wire       [5:0]    _zz_when_ArraySlice_l112_169;
  wire                when_ArraySlice_l112_169;
  wire                when_ArraySlice_l113_169;
  wire                when_ArraySlice_l118_169;
  wire                when_ArraySlice_l173_169;
  wire                when_ArraySlice_l165_170;
  wire                when_ArraySlice_l166_170;
  reg        [6:0]    _zz_when_ArraySlice_l173_170;
  wire       [5:0]    _zz_when_ArraySlice_l112_170;
  wire                when_ArraySlice_l112_170;
  wire                when_ArraySlice_l113_170;
  wire                when_ArraySlice_l118_170;
  wire                when_ArraySlice_l173_170;
  wire                when_ArraySlice_l165_171;
  wire                when_ArraySlice_l166_171;
  reg        [6:0]    _zz_when_ArraySlice_l173_171;
  wire       [5:0]    _zz_when_ArraySlice_l112_171;
  wire                when_ArraySlice_l112_171;
  wire                when_ArraySlice_l113_171;
  wire                when_ArraySlice_l118_171;
  wire                when_ArraySlice_l173_171;
  wire                when_ArraySlice_l165_172;
  wire                when_ArraySlice_l166_172;
  reg        [6:0]    _zz_when_ArraySlice_l173_172;
  wire       [5:0]    _zz_when_ArraySlice_l112_172;
  wire                when_ArraySlice_l112_172;
  wire                when_ArraySlice_l113_172;
  wire                when_ArraySlice_l118_172;
  wire                when_ArraySlice_l173_172;
  wire                when_ArraySlice_l165_173;
  wire                when_ArraySlice_l166_173;
  reg        [6:0]    _zz_when_ArraySlice_l173_173;
  wire       [5:0]    _zz_when_ArraySlice_l112_173;
  wire                when_ArraySlice_l112_173;
  wire                when_ArraySlice_l113_173;
  wire                when_ArraySlice_l118_173;
  wire                when_ArraySlice_l173_173;
  wire                when_ArraySlice_l165_174;
  wire                when_ArraySlice_l166_174;
  reg        [6:0]    _zz_when_ArraySlice_l173_174;
  wire       [5:0]    _zz_when_ArraySlice_l112_174;
  wire                when_ArraySlice_l112_174;
  wire                when_ArraySlice_l113_174;
  wire                when_ArraySlice_l118_174;
  wire                when_ArraySlice_l173_174;
  wire                when_ArraySlice_l165_175;
  wire                when_ArraySlice_l166_175;
  reg        [6:0]    _zz_when_ArraySlice_l173_175;
  wire       [5:0]    _zz_when_ArraySlice_l112_175;
  wire                when_ArraySlice_l112_175;
  wire                when_ArraySlice_l113_175;
  wire                when_ArraySlice_l118_175;
  wire                when_ArraySlice_l173_175;
  wire                when_ArraySlice_l444_6;
  wire                outputStreamArrayData_6_fire_5;
  wire                when_ArraySlice_l448_6;
  wire                when_ArraySlice_l434_6;
  wire                outputStreamArrayData_6_fire_6;
  wire                when_ArraySlice_l455_6;
  wire                when_ArraySlice_l373_7;
  wire                when_ArraySlice_l374_7;
  wire       [5:0]    _zz_outputStreamArrayData_7_valid;
  wire                _zz_io_pop_ready_7;
  wire       [63:0]   _zz_10;
  wire                when_ArraySlice_l379_7;
  wire                outputStreamArrayData_7_fire;
  wire                when_ArraySlice_l380_7;
  wire                when_ArraySlice_l381_7;
  wire                when_ArraySlice_l384_7;
  wire                outputStreamArrayData_7_fire_1;
  wire                when_ArraySlice_l389_7;
  wire                when_ArraySlice_l390_7;
  reg        [6:0]    _zz_when_ArraySlice_l392_7;
  wire       [5:0]    _zz_when_ArraySlice_l94_21;
  wire                when_ArraySlice_l94_21;
  wire                when_ArraySlice_l95_21;
  wire                when_ArraySlice_l99_21;
  wire                when_ArraySlice_l392_7;
  reg                 debug_0_22 /* verilator public */ ;
  reg                 debug_1_22 /* verilator public */ ;
  reg                 debug_2_22 /* verilator public */ ;
  reg                 debug_3_22 /* verilator public */ ;
  reg                 debug_4_22 /* verilator public */ ;
  reg                 debug_5_22 /* verilator public */ ;
  reg                 debug_6_22 /* verilator public */ ;
  reg                 debug_7_22 /* verilator public */ ;
  wire                when_ArraySlice_l165_176;
  wire                when_ArraySlice_l166_176;
  reg        [6:0]    _zz_when_ArraySlice_l173_176;
  wire       [5:0]    _zz_when_ArraySlice_l112_176;
  wire                when_ArraySlice_l112_176;
  wire                when_ArraySlice_l113_176;
  wire                when_ArraySlice_l118_176;
  wire                when_ArraySlice_l173_176;
  wire                when_ArraySlice_l165_177;
  wire                when_ArraySlice_l166_177;
  reg        [6:0]    _zz_when_ArraySlice_l173_177;
  wire       [5:0]    _zz_when_ArraySlice_l112_177;
  wire                when_ArraySlice_l112_177;
  wire                when_ArraySlice_l113_177;
  wire                when_ArraySlice_l118_177;
  wire                when_ArraySlice_l173_177;
  wire                when_ArraySlice_l165_178;
  wire                when_ArraySlice_l166_178;
  reg        [6:0]    _zz_when_ArraySlice_l173_178;
  wire       [5:0]    _zz_when_ArraySlice_l112_178;
  wire                when_ArraySlice_l112_178;
  wire                when_ArraySlice_l113_178;
  wire                when_ArraySlice_l118_178;
  wire                when_ArraySlice_l173_178;
  wire                when_ArraySlice_l165_179;
  wire                when_ArraySlice_l166_179;
  reg        [6:0]    _zz_when_ArraySlice_l173_179;
  wire       [5:0]    _zz_when_ArraySlice_l112_179;
  wire                when_ArraySlice_l112_179;
  wire                when_ArraySlice_l113_179;
  wire                when_ArraySlice_l118_179;
  wire                when_ArraySlice_l173_179;
  wire                when_ArraySlice_l165_180;
  wire                when_ArraySlice_l166_180;
  reg        [6:0]    _zz_when_ArraySlice_l173_180;
  wire       [5:0]    _zz_when_ArraySlice_l112_180;
  wire                when_ArraySlice_l112_180;
  wire                when_ArraySlice_l113_180;
  wire                when_ArraySlice_l118_180;
  wire                when_ArraySlice_l173_180;
  wire                when_ArraySlice_l165_181;
  wire                when_ArraySlice_l166_181;
  reg        [6:0]    _zz_when_ArraySlice_l173_181;
  wire       [5:0]    _zz_when_ArraySlice_l112_181;
  wire                when_ArraySlice_l112_181;
  wire                when_ArraySlice_l113_181;
  wire                when_ArraySlice_l118_181;
  wire                when_ArraySlice_l173_181;
  wire                when_ArraySlice_l165_182;
  wire                when_ArraySlice_l166_182;
  reg        [6:0]    _zz_when_ArraySlice_l173_182;
  wire       [5:0]    _zz_when_ArraySlice_l112_182;
  wire                when_ArraySlice_l112_182;
  wire                when_ArraySlice_l113_182;
  wire                when_ArraySlice_l118_182;
  wire                when_ArraySlice_l173_182;
  wire                when_ArraySlice_l165_183;
  wire                when_ArraySlice_l166_183;
  reg        [6:0]    _zz_when_ArraySlice_l173_183;
  wire       [5:0]    _zz_when_ArraySlice_l112_183;
  wire                when_ArraySlice_l112_183;
  wire                when_ArraySlice_l113_183;
  wire                when_ArraySlice_l118_183;
  wire                when_ArraySlice_l173_183;
  wire                when_ArraySlice_l398_7;
  wire                when_ArraySlice_l401_7;
  wire                when_ArraySlice_l405_7;
  wire                when_ArraySlice_l409_7;
  wire                outputStreamArrayData_7_fire_2;
  wire                when_ArraySlice_l410_7;
  reg        [6:0]    _zz_when_ArraySlice_l412_7;
  wire       [5:0]    _zz_when_ArraySlice_l94_22;
  wire                when_ArraySlice_l94_22;
  wire                when_ArraySlice_l95_22;
  wire                when_ArraySlice_l99_22;
  wire                when_ArraySlice_l412_7;
  reg                 debug_0_23 /* verilator public */ ;
  reg                 debug_1_23 /* verilator public */ ;
  reg                 debug_2_23 /* verilator public */ ;
  reg                 debug_3_23 /* verilator public */ ;
  reg                 debug_4_23 /* verilator public */ ;
  reg                 debug_5_23 /* verilator public */ ;
  reg                 debug_6_23 /* verilator public */ ;
  reg                 debug_7_23 /* verilator public */ ;
  wire                when_ArraySlice_l165_184;
  wire                when_ArraySlice_l166_184;
  reg        [6:0]    _zz_when_ArraySlice_l173_184;
  wire       [5:0]    _zz_when_ArraySlice_l112_184;
  wire                when_ArraySlice_l112_184;
  wire                when_ArraySlice_l113_184;
  wire                when_ArraySlice_l118_184;
  wire                when_ArraySlice_l173_184;
  wire                when_ArraySlice_l165_185;
  wire                when_ArraySlice_l166_185;
  reg        [6:0]    _zz_when_ArraySlice_l173_185;
  wire       [5:0]    _zz_when_ArraySlice_l112_185;
  wire                when_ArraySlice_l112_185;
  wire                when_ArraySlice_l113_185;
  wire                when_ArraySlice_l118_185;
  wire                when_ArraySlice_l173_185;
  wire                when_ArraySlice_l165_186;
  wire                when_ArraySlice_l166_186;
  reg        [6:0]    _zz_when_ArraySlice_l173_186;
  wire       [5:0]    _zz_when_ArraySlice_l112_186;
  wire                when_ArraySlice_l112_186;
  wire                when_ArraySlice_l113_186;
  wire                when_ArraySlice_l118_186;
  wire                when_ArraySlice_l173_186;
  wire                when_ArraySlice_l165_187;
  wire                when_ArraySlice_l166_187;
  reg        [6:0]    _zz_when_ArraySlice_l173_187;
  wire       [5:0]    _zz_when_ArraySlice_l112_187;
  wire                when_ArraySlice_l112_187;
  wire                when_ArraySlice_l113_187;
  wire                when_ArraySlice_l118_187;
  wire                when_ArraySlice_l173_187;
  wire                when_ArraySlice_l165_188;
  wire                when_ArraySlice_l166_188;
  reg        [6:0]    _zz_when_ArraySlice_l173_188;
  wire       [5:0]    _zz_when_ArraySlice_l112_188;
  wire                when_ArraySlice_l112_188;
  wire                when_ArraySlice_l113_188;
  wire                when_ArraySlice_l118_188;
  wire                when_ArraySlice_l173_188;
  wire                when_ArraySlice_l165_189;
  wire                when_ArraySlice_l166_189;
  reg        [6:0]    _zz_when_ArraySlice_l173_189;
  wire       [5:0]    _zz_when_ArraySlice_l112_189;
  wire                when_ArraySlice_l112_189;
  wire                when_ArraySlice_l113_189;
  wire                when_ArraySlice_l118_189;
  wire                when_ArraySlice_l173_189;
  wire                when_ArraySlice_l165_190;
  wire                when_ArraySlice_l166_190;
  reg        [6:0]    _zz_when_ArraySlice_l173_190;
  wire       [5:0]    _zz_when_ArraySlice_l112_190;
  wire                when_ArraySlice_l112_190;
  wire                when_ArraySlice_l113_190;
  wire                when_ArraySlice_l118_190;
  wire                when_ArraySlice_l173_190;
  wire                when_ArraySlice_l165_191;
  wire                when_ArraySlice_l166_191;
  reg        [6:0]    _zz_when_ArraySlice_l173_191;
  wire       [5:0]    _zz_when_ArraySlice_l112_191;
  wire                when_ArraySlice_l112_191;
  wire                when_ArraySlice_l113_191;
  wire                when_ArraySlice_l118_191;
  wire                when_ArraySlice_l173_191;
  wire                when_ArraySlice_l418_7;
  wire                when_ArraySlice_l421_7;
  wire                outputStreamArrayData_7_fire_3;
  wire                when_ArraySlice_l425_7;
  wire                outputStreamArrayData_7_fire_4;
  wire                when_ArraySlice_l436_7;
  reg        [6:0]    _zz_when_ArraySlice_l437_7;
  wire       [5:0]    _zz_when_ArraySlice_l94_23;
  wire                when_ArraySlice_l94_23;
  wire                when_ArraySlice_l95_23;
  wire                when_ArraySlice_l99_23;
  wire                when_ArraySlice_l437_7;
  reg                 debug_0_24 /* verilator public */ ;
  reg                 debug_1_24 /* verilator public */ ;
  reg                 debug_2_24 /* verilator public */ ;
  reg                 debug_3_24 /* verilator public */ ;
  reg                 debug_4_24 /* verilator public */ ;
  reg                 debug_5_24 /* verilator public */ ;
  reg                 debug_6_24 /* verilator public */ ;
  reg                 debug_7_24 /* verilator public */ ;
  wire                when_ArraySlice_l165_192;
  wire                when_ArraySlice_l166_192;
  reg        [6:0]    _zz_when_ArraySlice_l173_192;
  wire       [5:0]    _zz_when_ArraySlice_l112_192;
  wire                when_ArraySlice_l112_192;
  wire                when_ArraySlice_l113_192;
  wire                when_ArraySlice_l118_192;
  wire                when_ArraySlice_l173_192;
  wire                when_ArraySlice_l165_193;
  wire                when_ArraySlice_l166_193;
  reg        [6:0]    _zz_when_ArraySlice_l173_193;
  wire       [5:0]    _zz_when_ArraySlice_l112_193;
  wire                when_ArraySlice_l112_193;
  wire                when_ArraySlice_l113_193;
  wire                when_ArraySlice_l118_193;
  wire                when_ArraySlice_l173_193;
  wire                when_ArraySlice_l165_194;
  wire                when_ArraySlice_l166_194;
  reg        [6:0]    _zz_when_ArraySlice_l173_194;
  wire       [5:0]    _zz_when_ArraySlice_l112_194;
  wire                when_ArraySlice_l112_194;
  wire                when_ArraySlice_l113_194;
  wire                when_ArraySlice_l118_194;
  wire                when_ArraySlice_l173_194;
  wire                when_ArraySlice_l165_195;
  wire                when_ArraySlice_l166_195;
  reg        [6:0]    _zz_when_ArraySlice_l173_195;
  wire       [5:0]    _zz_when_ArraySlice_l112_195;
  wire                when_ArraySlice_l112_195;
  wire                when_ArraySlice_l113_195;
  wire                when_ArraySlice_l118_195;
  wire                when_ArraySlice_l173_195;
  wire                when_ArraySlice_l165_196;
  wire                when_ArraySlice_l166_196;
  reg        [6:0]    _zz_when_ArraySlice_l173_196;
  wire       [5:0]    _zz_when_ArraySlice_l112_196;
  wire                when_ArraySlice_l112_196;
  wire                when_ArraySlice_l113_196;
  wire                when_ArraySlice_l118_196;
  wire                when_ArraySlice_l173_196;
  wire                when_ArraySlice_l165_197;
  wire                when_ArraySlice_l166_197;
  reg        [6:0]    _zz_when_ArraySlice_l173_197;
  wire       [5:0]    _zz_when_ArraySlice_l112_197;
  wire                when_ArraySlice_l112_197;
  wire                when_ArraySlice_l113_197;
  wire                when_ArraySlice_l118_197;
  wire                when_ArraySlice_l173_197;
  wire                when_ArraySlice_l165_198;
  wire                when_ArraySlice_l166_198;
  reg        [6:0]    _zz_when_ArraySlice_l173_198;
  wire       [5:0]    _zz_when_ArraySlice_l112_198;
  wire                when_ArraySlice_l112_198;
  wire                when_ArraySlice_l113_198;
  wire                when_ArraySlice_l118_198;
  wire                when_ArraySlice_l173_198;
  wire                when_ArraySlice_l165_199;
  wire                when_ArraySlice_l166_199;
  reg        [6:0]    _zz_when_ArraySlice_l173_199;
  wire       [5:0]    _zz_when_ArraySlice_l112_199;
  wire                when_ArraySlice_l112_199;
  wire                when_ArraySlice_l113_199;
  wire                when_ArraySlice_l118_199;
  wire                when_ArraySlice_l173_199;
  wire                when_ArraySlice_l444_7;
  wire                outputStreamArrayData_7_fire_5;
  wire                when_ArraySlice_l448_7;
  wire                when_ArraySlice_l434_7;
  wire                outputStreamArrayData_7_fire_6;
  wire                when_ArraySlice_l455_7;
  reg                 debug_0_25 /* verilator public */ ;
  reg                 debug_1_25 /* verilator public */ ;
  reg                 debug_2_25 /* verilator public */ ;
  reg                 debug_3_25 /* verilator public */ ;
  reg                 debug_4_25 /* verilator public */ ;
  reg                 debug_5_25 /* verilator public */ ;
  reg                 debug_6_25 /* verilator public */ ;
  reg                 debug_7_25 /* verilator public */ ;
  wire                when_ArraySlice_l165_200;
  wire                when_ArraySlice_l166_200;
  reg        [6:0]    _zz_when_ArraySlice_l173_200;
  wire       [5:0]    _zz_when_ArraySlice_l112_200;
  wire                when_ArraySlice_l112_200;
  wire                when_ArraySlice_l113_200;
  wire                when_ArraySlice_l118_200;
  wire                when_ArraySlice_l173_200;
  wire                when_ArraySlice_l165_201;
  wire                when_ArraySlice_l166_201;
  reg        [6:0]    _zz_when_ArraySlice_l173_201;
  wire       [5:0]    _zz_when_ArraySlice_l112_201;
  wire                when_ArraySlice_l112_201;
  wire                when_ArraySlice_l113_201;
  wire                when_ArraySlice_l118_201;
  wire                when_ArraySlice_l173_201;
  wire                when_ArraySlice_l165_202;
  wire                when_ArraySlice_l166_202;
  reg        [6:0]    _zz_when_ArraySlice_l173_202;
  wire       [5:0]    _zz_when_ArraySlice_l112_202;
  wire                when_ArraySlice_l112_202;
  wire                when_ArraySlice_l113_202;
  wire                when_ArraySlice_l118_202;
  wire                when_ArraySlice_l173_202;
  wire                when_ArraySlice_l165_203;
  wire                when_ArraySlice_l166_203;
  reg        [6:0]    _zz_when_ArraySlice_l173_203;
  wire       [5:0]    _zz_when_ArraySlice_l112_203;
  wire                when_ArraySlice_l112_203;
  wire                when_ArraySlice_l113_203;
  wire                when_ArraySlice_l118_203;
  wire                when_ArraySlice_l173_203;
  wire                when_ArraySlice_l165_204;
  wire                when_ArraySlice_l166_204;
  reg        [6:0]    _zz_when_ArraySlice_l173_204;
  wire       [5:0]    _zz_when_ArraySlice_l112_204;
  wire                when_ArraySlice_l112_204;
  wire                when_ArraySlice_l113_204;
  wire                when_ArraySlice_l118_204;
  wire                when_ArraySlice_l173_204;
  wire                when_ArraySlice_l165_205;
  wire                when_ArraySlice_l166_205;
  reg        [6:0]    _zz_when_ArraySlice_l173_205;
  wire       [5:0]    _zz_when_ArraySlice_l112_205;
  wire                when_ArraySlice_l112_205;
  wire                when_ArraySlice_l113_205;
  wire                when_ArraySlice_l118_205;
  wire                when_ArraySlice_l173_205;
  wire                when_ArraySlice_l165_206;
  wire                when_ArraySlice_l166_206;
  reg        [6:0]    _zz_when_ArraySlice_l173_206;
  wire       [5:0]    _zz_when_ArraySlice_l112_206;
  wire                when_ArraySlice_l112_206;
  wire                when_ArraySlice_l113_206;
  wire                when_ArraySlice_l118_206;
  wire                when_ArraySlice_l173_206;
  wire                when_ArraySlice_l165_207;
  wire                when_ArraySlice_l166_207;
  reg        [6:0]    _zz_when_ArraySlice_l173_207;
  wire       [5:0]    _zz_when_ArraySlice_l112_207;
  wire                when_ArraySlice_l112_207;
  wire                when_ArraySlice_l113_207;
  wire                when_ArraySlice_l118_207;
  wire                when_ArraySlice_l173_207;
  wire                when_ArraySlice_l465;
  wire                when_ArraySlice_l468;
  wire                when_ArraySlice_l468_1;
  wire                when_ArraySlice_l468_2;
  wire                when_ArraySlice_l468_3;
  wire                when_ArraySlice_l468_4;
  wire                when_ArraySlice_l468_5;
  wire                when_ArraySlice_l468_6;
  wire                when_ArraySlice_l468_7;
  wire                when_ArraySlice_l240;
  wire                when_ArraySlice_l241;
  wire       [5:0]    _zz_outputStreamArrayData_0_valid_1;
  wire                _zz_io_pop_ready_8;
  wire       [63:0]   _zz_11;
  wire                when_ArraySlice_l246;
  wire                outputStreamArrayData_0_fire_7;
  wire                when_ArraySlice_l247;
  wire                when_ArraySlice_l248;
  wire                when_ArraySlice_l251;
  wire                outputStreamArrayData_0_fire_8;
  wire                when_ArraySlice_l256;
  wire                when_ArraySlice_l257;
  reg        [6:0]    _zz_when_ArraySlice_l259;
  wire       [5:0]    _zz_when_ArraySlice_l94_24;
  wire                when_ArraySlice_l94_24;
  wire                when_ArraySlice_l95_24;
  wire                when_ArraySlice_l99_24;
  wire                when_ArraySlice_l259;
  reg                 debug_0_26 /* verilator public */ ;
  reg                 debug_1_26 /* verilator public */ ;
  reg                 debug_2_26 /* verilator public */ ;
  reg                 debug_3_26 /* verilator public */ ;
  reg                 debug_4_26 /* verilator public */ ;
  reg                 debug_5_26 /* verilator public */ ;
  reg                 debug_6_26 /* verilator public */ ;
  reg                 debug_7_26 /* verilator public */ ;
  wire                when_ArraySlice_l165_208;
  wire                when_ArraySlice_l166_208;
  reg        [6:0]    _zz_when_ArraySlice_l173_208;
  wire       [5:0]    _zz_when_ArraySlice_l112_208;
  wire                when_ArraySlice_l112_208;
  wire                when_ArraySlice_l113_208;
  wire                when_ArraySlice_l118_208;
  wire                when_ArraySlice_l173_208;
  wire                when_ArraySlice_l165_209;
  wire                when_ArraySlice_l166_209;
  reg        [6:0]    _zz_when_ArraySlice_l173_209;
  wire       [5:0]    _zz_when_ArraySlice_l112_209;
  wire                when_ArraySlice_l112_209;
  wire                when_ArraySlice_l113_209;
  wire                when_ArraySlice_l118_209;
  wire                when_ArraySlice_l173_209;
  wire                when_ArraySlice_l165_210;
  wire                when_ArraySlice_l166_210;
  reg        [6:0]    _zz_when_ArraySlice_l173_210;
  wire       [5:0]    _zz_when_ArraySlice_l112_210;
  wire                when_ArraySlice_l112_210;
  wire                when_ArraySlice_l113_210;
  wire                when_ArraySlice_l118_210;
  wire                when_ArraySlice_l173_210;
  wire                when_ArraySlice_l165_211;
  wire                when_ArraySlice_l166_211;
  reg        [6:0]    _zz_when_ArraySlice_l173_211;
  wire       [5:0]    _zz_when_ArraySlice_l112_211;
  wire                when_ArraySlice_l112_211;
  wire                when_ArraySlice_l113_211;
  wire                when_ArraySlice_l118_211;
  wire                when_ArraySlice_l173_211;
  wire                when_ArraySlice_l165_212;
  wire                when_ArraySlice_l166_212;
  reg        [6:0]    _zz_when_ArraySlice_l173_212;
  wire       [5:0]    _zz_when_ArraySlice_l112_212;
  wire                when_ArraySlice_l112_212;
  wire                when_ArraySlice_l113_212;
  wire                when_ArraySlice_l118_212;
  wire                when_ArraySlice_l173_212;
  wire                when_ArraySlice_l165_213;
  wire                when_ArraySlice_l166_213;
  reg        [6:0]    _zz_when_ArraySlice_l173_213;
  wire       [5:0]    _zz_when_ArraySlice_l112_213;
  wire                when_ArraySlice_l112_213;
  wire                when_ArraySlice_l113_213;
  wire                when_ArraySlice_l118_213;
  wire                when_ArraySlice_l173_213;
  wire                when_ArraySlice_l165_214;
  wire                when_ArraySlice_l166_214;
  reg        [6:0]    _zz_when_ArraySlice_l173_214;
  wire       [5:0]    _zz_when_ArraySlice_l112_214;
  wire                when_ArraySlice_l112_214;
  wire                when_ArraySlice_l113_214;
  wire                when_ArraySlice_l118_214;
  wire                when_ArraySlice_l173_214;
  wire                when_ArraySlice_l165_215;
  wire                when_ArraySlice_l166_215;
  reg        [6:0]    _zz_when_ArraySlice_l173_215;
  wire       [5:0]    _zz_when_ArraySlice_l112_215;
  wire                when_ArraySlice_l112_215;
  wire                when_ArraySlice_l113_215;
  wire                when_ArraySlice_l118_215;
  wire                when_ArraySlice_l173_215;
  wire                when_ArraySlice_l265;
  wire                when_ArraySlice_l268;
  wire                when_ArraySlice_l272;
  wire                when_ArraySlice_l276;
  wire                outputStreamArrayData_0_fire_9;
  wire                when_ArraySlice_l277;
  reg        [6:0]    _zz_when_ArraySlice_l279;
  wire       [5:0]    _zz_when_ArraySlice_l94_25;
  wire                when_ArraySlice_l94_25;
  wire                when_ArraySlice_l95_25;
  wire                when_ArraySlice_l99_25;
  wire                when_ArraySlice_l279;
  reg                 debug_0_27 /* verilator public */ ;
  reg                 debug_1_27 /* verilator public */ ;
  reg                 debug_2_27 /* verilator public */ ;
  reg                 debug_3_27 /* verilator public */ ;
  reg                 debug_4_27 /* verilator public */ ;
  reg                 debug_5_27 /* verilator public */ ;
  reg                 debug_6_27 /* verilator public */ ;
  reg                 debug_7_27 /* verilator public */ ;
  wire                when_ArraySlice_l165_216;
  wire                when_ArraySlice_l166_216;
  reg        [6:0]    _zz_when_ArraySlice_l173_216;
  wire       [5:0]    _zz_when_ArraySlice_l112_216;
  wire                when_ArraySlice_l112_216;
  wire                when_ArraySlice_l113_216;
  wire                when_ArraySlice_l118_216;
  wire                when_ArraySlice_l173_216;
  wire                when_ArraySlice_l165_217;
  wire                when_ArraySlice_l166_217;
  reg        [6:0]    _zz_when_ArraySlice_l173_217;
  wire       [5:0]    _zz_when_ArraySlice_l112_217;
  wire                when_ArraySlice_l112_217;
  wire                when_ArraySlice_l113_217;
  wire                when_ArraySlice_l118_217;
  wire                when_ArraySlice_l173_217;
  wire                when_ArraySlice_l165_218;
  wire                when_ArraySlice_l166_218;
  reg        [6:0]    _zz_when_ArraySlice_l173_218;
  wire       [5:0]    _zz_when_ArraySlice_l112_218;
  wire                when_ArraySlice_l112_218;
  wire                when_ArraySlice_l113_218;
  wire                when_ArraySlice_l118_218;
  wire                when_ArraySlice_l173_218;
  wire                when_ArraySlice_l165_219;
  wire                when_ArraySlice_l166_219;
  reg        [6:0]    _zz_when_ArraySlice_l173_219;
  wire       [5:0]    _zz_when_ArraySlice_l112_219;
  wire                when_ArraySlice_l112_219;
  wire                when_ArraySlice_l113_219;
  wire                when_ArraySlice_l118_219;
  wire                when_ArraySlice_l173_219;
  wire                when_ArraySlice_l165_220;
  wire                when_ArraySlice_l166_220;
  reg        [6:0]    _zz_when_ArraySlice_l173_220;
  wire       [5:0]    _zz_when_ArraySlice_l112_220;
  wire                when_ArraySlice_l112_220;
  wire                when_ArraySlice_l113_220;
  wire                when_ArraySlice_l118_220;
  wire                when_ArraySlice_l173_220;
  wire                when_ArraySlice_l165_221;
  wire                when_ArraySlice_l166_221;
  reg        [6:0]    _zz_when_ArraySlice_l173_221;
  wire       [5:0]    _zz_when_ArraySlice_l112_221;
  wire                when_ArraySlice_l112_221;
  wire                when_ArraySlice_l113_221;
  wire                when_ArraySlice_l118_221;
  wire                when_ArraySlice_l173_221;
  wire                when_ArraySlice_l165_222;
  wire                when_ArraySlice_l166_222;
  reg        [6:0]    _zz_when_ArraySlice_l173_222;
  wire       [5:0]    _zz_when_ArraySlice_l112_222;
  wire                when_ArraySlice_l112_222;
  wire                when_ArraySlice_l113_222;
  wire                when_ArraySlice_l118_222;
  wire                when_ArraySlice_l173_222;
  wire                when_ArraySlice_l165_223;
  wire                when_ArraySlice_l166_223;
  reg        [6:0]    _zz_when_ArraySlice_l173_223;
  wire       [5:0]    _zz_when_ArraySlice_l112_223;
  wire                when_ArraySlice_l112_223;
  wire                when_ArraySlice_l113_223;
  wire                when_ArraySlice_l118_223;
  wire                when_ArraySlice_l173_223;
  wire                when_ArraySlice_l285;
  wire                when_ArraySlice_l288;
  wire                outputStreamArrayData_0_fire_10;
  wire                when_ArraySlice_l292;
  wire                outputStreamArrayData_0_fire_11;
  wire                when_ArraySlice_l303;
  reg        [6:0]    _zz_when_ArraySlice_l304;
  wire       [5:0]    _zz_when_ArraySlice_l94_26;
  wire                when_ArraySlice_l94_26;
  wire                when_ArraySlice_l95_26;
  wire                when_ArraySlice_l99_26;
  wire                when_ArraySlice_l304;
  reg                 debug_0_28 /* verilator public */ ;
  reg                 debug_1_28 /* verilator public */ ;
  reg                 debug_2_28 /* verilator public */ ;
  reg                 debug_3_28 /* verilator public */ ;
  reg                 debug_4_28 /* verilator public */ ;
  reg                 debug_5_28 /* verilator public */ ;
  reg                 debug_6_28 /* verilator public */ ;
  reg                 debug_7_28 /* verilator public */ ;
  wire                when_ArraySlice_l165_224;
  wire                when_ArraySlice_l166_224;
  reg        [6:0]    _zz_when_ArraySlice_l173_224;
  wire       [5:0]    _zz_when_ArraySlice_l112_224;
  wire                when_ArraySlice_l112_224;
  wire                when_ArraySlice_l113_224;
  wire                when_ArraySlice_l118_224;
  wire                when_ArraySlice_l173_224;
  wire                when_ArraySlice_l165_225;
  wire                when_ArraySlice_l166_225;
  reg        [6:0]    _zz_when_ArraySlice_l173_225;
  wire       [5:0]    _zz_when_ArraySlice_l112_225;
  wire                when_ArraySlice_l112_225;
  wire                when_ArraySlice_l113_225;
  wire                when_ArraySlice_l118_225;
  wire                when_ArraySlice_l173_225;
  wire                when_ArraySlice_l165_226;
  wire                when_ArraySlice_l166_226;
  reg        [6:0]    _zz_when_ArraySlice_l173_226;
  wire       [5:0]    _zz_when_ArraySlice_l112_226;
  wire                when_ArraySlice_l112_226;
  wire                when_ArraySlice_l113_226;
  wire                when_ArraySlice_l118_226;
  wire                when_ArraySlice_l173_226;
  wire                when_ArraySlice_l165_227;
  wire                when_ArraySlice_l166_227;
  reg        [6:0]    _zz_when_ArraySlice_l173_227;
  wire       [5:0]    _zz_when_ArraySlice_l112_227;
  wire                when_ArraySlice_l112_227;
  wire                when_ArraySlice_l113_227;
  wire                when_ArraySlice_l118_227;
  wire                when_ArraySlice_l173_227;
  wire                when_ArraySlice_l165_228;
  wire                when_ArraySlice_l166_228;
  reg        [6:0]    _zz_when_ArraySlice_l173_228;
  wire       [5:0]    _zz_when_ArraySlice_l112_228;
  wire                when_ArraySlice_l112_228;
  wire                when_ArraySlice_l113_228;
  wire                when_ArraySlice_l118_228;
  wire                when_ArraySlice_l173_228;
  wire                when_ArraySlice_l165_229;
  wire                when_ArraySlice_l166_229;
  reg        [6:0]    _zz_when_ArraySlice_l173_229;
  wire       [5:0]    _zz_when_ArraySlice_l112_229;
  wire                when_ArraySlice_l112_229;
  wire                when_ArraySlice_l113_229;
  wire                when_ArraySlice_l118_229;
  wire                when_ArraySlice_l173_229;
  wire                when_ArraySlice_l165_230;
  wire                when_ArraySlice_l166_230;
  reg        [6:0]    _zz_when_ArraySlice_l173_230;
  wire       [5:0]    _zz_when_ArraySlice_l112_230;
  wire                when_ArraySlice_l112_230;
  wire                when_ArraySlice_l113_230;
  wire                when_ArraySlice_l118_230;
  wire                when_ArraySlice_l173_230;
  wire                when_ArraySlice_l165_231;
  wire                when_ArraySlice_l166_231;
  reg        [6:0]    _zz_when_ArraySlice_l173_231;
  wire       [5:0]    _zz_when_ArraySlice_l112_231;
  wire                when_ArraySlice_l112_231;
  wire                when_ArraySlice_l113_231;
  wire                when_ArraySlice_l118_231;
  wire                when_ArraySlice_l173_231;
  wire                when_ArraySlice_l311;
  wire                outputStreamArrayData_0_fire_12;
  wire                when_ArraySlice_l315;
  wire                when_ArraySlice_l301;
  wire                outputStreamArrayData_0_fire_13;
  wire                when_ArraySlice_l322;
  wire                when_ArraySlice_l240_1;
  wire                when_ArraySlice_l241_1;
  wire       [5:0]    _zz_outputStreamArrayData_1_valid_1;
  wire                _zz_io_pop_ready_9;
  wire       [63:0]   _zz_12;
  wire                when_ArraySlice_l246_1;
  wire                outputStreamArrayData_1_fire_7;
  wire                when_ArraySlice_l247_1;
  wire                when_ArraySlice_l248_1;
  wire                when_ArraySlice_l251_1;
  wire                outputStreamArrayData_1_fire_8;
  wire                when_ArraySlice_l256_1;
  wire                when_ArraySlice_l257_1;
  reg        [6:0]    _zz_when_ArraySlice_l259_1;
  wire       [5:0]    _zz_when_ArraySlice_l94_27;
  wire                when_ArraySlice_l94_27;
  wire                when_ArraySlice_l95_27;
  wire                when_ArraySlice_l99_27;
  wire                when_ArraySlice_l259_1;
  reg                 debug_0_29 /* verilator public */ ;
  reg                 debug_1_29 /* verilator public */ ;
  reg                 debug_2_29 /* verilator public */ ;
  reg                 debug_3_29 /* verilator public */ ;
  reg                 debug_4_29 /* verilator public */ ;
  reg                 debug_5_29 /* verilator public */ ;
  reg                 debug_6_29 /* verilator public */ ;
  reg                 debug_7_29 /* verilator public */ ;
  wire                when_ArraySlice_l165_232;
  wire                when_ArraySlice_l166_232;
  reg        [6:0]    _zz_when_ArraySlice_l173_232;
  wire       [5:0]    _zz_when_ArraySlice_l112_232;
  wire                when_ArraySlice_l112_232;
  wire                when_ArraySlice_l113_232;
  wire                when_ArraySlice_l118_232;
  wire                when_ArraySlice_l173_232;
  wire                when_ArraySlice_l165_233;
  wire                when_ArraySlice_l166_233;
  reg        [6:0]    _zz_when_ArraySlice_l173_233;
  wire       [5:0]    _zz_when_ArraySlice_l112_233;
  wire                when_ArraySlice_l112_233;
  wire                when_ArraySlice_l113_233;
  wire                when_ArraySlice_l118_233;
  wire                when_ArraySlice_l173_233;
  wire                when_ArraySlice_l165_234;
  wire                when_ArraySlice_l166_234;
  reg        [6:0]    _zz_when_ArraySlice_l173_234;
  wire       [5:0]    _zz_when_ArraySlice_l112_234;
  wire                when_ArraySlice_l112_234;
  wire                when_ArraySlice_l113_234;
  wire                when_ArraySlice_l118_234;
  wire                when_ArraySlice_l173_234;
  wire                when_ArraySlice_l165_235;
  wire                when_ArraySlice_l166_235;
  reg        [6:0]    _zz_when_ArraySlice_l173_235;
  wire       [5:0]    _zz_when_ArraySlice_l112_235;
  wire                when_ArraySlice_l112_235;
  wire                when_ArraySlice_l113_235;
  wire                when_ArraySlice_l118_235;
  wire                when_ArraySlice_l173_235;
  wire                when_ArraySlice_l165_236;
  wire                when_ArraySlice_l166_236;
  reg        [6:0]    _zz_when_ArraySlice_l173_236;
  wire       [5:0]    _zz_when_ArraySlice_l112_236;
  wire                when_ArraySlice_l112_236;
  wire                when_ArraySlice_l113_236;
  wire                when_ArraySlice_l118_236;
  wire                when_ArraySlice_l173_236;
  wire                when_ArraySlice_l165_237;
  wire                when_ArraySlice_l166_237;
  reg        [6:0]    _zz_when_ArraySlice_l173_237;
  wire       [5:0]    _zz_when_ArraySlice_l112_237;
  wire                when_ArraySlice_l112_237;
  wire                when_ArraySlice_l113_237;
  wire                when_ArraySlice_l118_237;
  wire                when_ArraySlice_l173_237;
  wire                when_ArraySlice_l165_238;
  wire                when_ArraySlice_l166_238;
  reg        [6:0]    _zz_when_ArraySlice_l173_238;
  wire       [5:0]    _zz_when_ArraySlice_l112_238;
  wire                when_ArraySlice_l112_238;
  wire                when_ArraySlice_l113_238;
  wire                when_ArraySlice_l118_238;
  wire                when_ArraySlice_l173_238;
  wire                when_ArraySlice_l165_239;
  wire                when_ArraySlice_l166_239;
  reg        [6:0]    _zz_when_ArraySlice_l173_239;
  wire       [5:0]    _zz_when_ArraySlice_l112_239;
  wire                when_ArraySlice_l112_239;
  wire                when_ArraySlice_l113_239;
  wire                when_ArraySlice_l118_239;
  wire                when_ArraySlice_l173_239;
  wire                when_ArraySlice_l265_1;
  wire                when_ArraySlice_l268_1;
  wire                when_ArraySlice_l272_1;
  wire                when_ArraySlice_l276_1;
  wire                outputStreamArrayData_1_fire_9;
  wire                when_ArraySlice_l277_1;
  reg        [6:0]    _zz_when_ArraySlice_l279_1;
  wire       [5:0]    _zz_when_ArraySlice_l94_28;
  wire                when_ArraySlice_l94_28;
  wire                when_ArraySlice_l95_28;
  wire                when_ArraySlice_l99_28;
  wire                when_ArraySlice_l279_1;
  reg                 debug_0_30 /* verilator public */ ;
  reg                 debug_1_30 /* verilator public */ ;
  reg                 debug_2_30 /* verilator public */ ;
  reg                 debug_3_30 /* verilator public */ ;
  reg                 debug_4_30 /* verilator public */ ;
  reg                 debug_5_30 /* verilator public */ ;
  reg                 debug_6_30 /* verilator public */ ;
  reg                 debug_7_30 /* verilator public */ ;
  wire                when_ArraySlice_l165_240;
  wire                when_ArraySlice_l166_240;
  reg        [6:0]    _zz_when_ArraySlice_l173_240;
  wire       [5:0]    _zz_when_ArraySlice_l112_240;
  wire                when_ArraySlice_l112_240;
  wire                when_ArraySlice_l113_240;
  wire                when_ArraySlice_l118_240;
  wire                when_ArraySlice_l173_240;
  wire                when_ArraySlice_l165_241;
  wire                when_ArraySlice_l166_241;
  reg        [6:0]    _zz_when_ArraySlice_l173_241;
  wire       [5:0]    _zz_when_ArraySlice_l112_241;
  wire                when_ArraySlice_l112_241;
  wire                when_ArraySlice_l113_241;
  wire                when_ArraySlice_l118_241;
  wire                when_ArraySlice_l173_241;
  wire                when_ArraySlice_l165_242;
  wire                when_ArraySlice_l166_242;
  reg        [6:0]    _zz_when_ArraySlice_l173_242;
  wire       [5:0]    _zz_when_ArraySlice_l112_242;
  wire                when_ArraySlice_l112_242;
  wire                when_ArraySlice_l113_242;
  wire                when_ArraySlice_l118_242;
  wire                when_ArraySlice_l173_242;
  wire                when_ArraySlice_l165_243;
  wire                when_ArraySlice_l166_243;
  reg        [6:0]    _zz_when_ArraySlice_l173_243;
  wire       [5:0]    _zz_when_ArraySlice_l112_243;
  wire                when_ArraySlice_l112_243;
  wire                when_ArraySlice_l113_243;
  wire                when_ArraySlice_l118_243;
  wire                when_ArraySlice_l173_243;
  wire                when_ArraySlice_l165_244;
  wire                when_ArraySlice_l166_244;
  reg        [6:0]    _zz_when_ArraySlice_l173_244;
  wire       [5:0]    _zz_when_ArraySlice_l112_244;
  wire                when_ArraySlice_l112_244;
  wire                when_ArraySlice_l113_244;
  wire                when_ArraySlice_l118_244;
  wire                when_ArraySlice_l173_244;
  wire                when_ArraySlice_l165_245;
  wire                when_ArraySlice_l166_245;
  reg        [6:0]    _zz_when_ArraySlice_l173_245;
  wire       [5:0]    _zz_when_ArraySlice_l112_245;
  wire                when_ArraySlice_l112_245;
  wire                when_ArraySlice_l113_245;
  wire                when_ArraySlice_l118_245;
  wire                when_ArraySlice_l173_245;
  wire                when_ArraySlice_l165_246;
  wire                when_ArraySlice_l166_246;
  reg        [6:0]    _zz_when_ArraySlice_l173_246;
  wire       [5:0]    _zz_when_ArraySlice_l112_246;
  wire                when_ArraySlice_l112_246;
  wire                when_ArraySlice_l113_246;
  wire                when_ArraySlice_l118_246;
  wire                when_ArraySlice_l173_246;
  wire                when_ArraySlice_l165_247;
  wire                when_ArraySlice_l166_247;
  reg        [6:0]    _zz_when_ArraySlice_l173_247;
  wire       [5:0]    _zz_when_ArraySlice_l112_247;
  wire                when_ArraySlice_l112_247;
  wire                when_ArraySlice_l113_247;
  wire                when_ArraySlice_l118_247;
  wire                when_ArraySlice_l173_247;
  wire                when_ArraySlice_l285_1;
  wire                when_ArraySlice_l288_1;
  wire                outputStreamArrayData_1_fire_10;
  wire                when_ArraySlice_l292_1;
  wire                outputStreamArrayData_1_fire_11;
  wire                when_ArraySlice_l303_1;
  reg        [6:0]    _zz_when_ArraySlice_l304_1;
  wire       [5:0]    _zz_when_ArraySlice_l94_29;
  wire                when_ArraySlice_l94_29;
  wire                when_ArraySlice_l95_29;
  wire                when_ArraySlice_l99_29;
  wire                when_ArraySlice_l304_1;
  reg                 debug_0_31 /* verilator public */ ;
  reg                 debug_1_31 /* verilator public */ ;
  reg                 debug_2_31 /* verilator public */ ;
  reg                 debug_3_31 /* verilator public */ ;
  reg                 debug_4_31 /* verilator public */ ;
  reg                 debug_5_31 /* verilator public */ ;
  reg                 debug_6_31 /* verilator public */ ;
  reg                 debug_7_31 /* verilator public */ ;
  wire                when_ArraySlice_l165_248;
  wire                when_ArraySlice_l166_248;
  reg        [6:0]    _zz_when_ArraySlice_l173_248;
  wire       [5:0]    _zz_when_ArraySlice_l112_248;
  wire                when_ArraySlice_l112_248;
  wire                when_ArraySlice_l113_248;
  wire                when_ArraySlice_l118_248;
  wire                when_ArraySlice_l173_248;
  wire                when_ArraySlice_l165_249;
  wire                when_ArraySlice_l166_249;
  reg        [6:0]    _zz_when_ArraySlice_l173_249;
  wire       [5:0]    _zz_when_ArraySlice_l112_249;
  wire                when_ArraySlice_l112_249;
  wire                when_ArraySlice_l113_249;
  wire                when_ArraySlice_l118_249;
  wire                when_ArraySlice_l173_249;
  wire                when_ArraySlice_l165_250;
  wire                when_ArraySlice_l166_250;
  reg        [6:0]    _zz_when_ArraySlice_l173_250;
  wire       [5:0]    _zz_when_ArraySlice_l112_250;
  wire                when_ArraySlice_l112_250;
  wire                when_ArraySlice_l113_250;
  wire                when_ArraySlice_l118_250;
  wire                when_ArraySlice_l173_250;
  wire                when_ArraySlice_l165_251;
  wire                when_ArraySlice_l166_251;
  reg        [6:0]    _zz_when_ArraySlice_l173_251;
  wire       [5:0]    _zz_when_ArraySlice_l112_251;
  wire                when_ArraySlice_l112_251;
  wire                when_ArraySlice_l113_251;
  wire                when_ArraySlice_l118_251;
  wire                when_ArraySlice_l173_251;
  wire                when_ArraySlice_l165_252;
  wire                when_ArraySlice_l166_252;
  reg        [6:0]    _zz_when_ArraySlice_l173_252;
  wire       [5:0]    _zz_when_ArraySlice_l112_252;
  wire                when_ArraySlice_l112_252;
  wire                when_ArraySlice_l113_252;
  wire                when_ArraySlice_l118_252;
  wire                when_ArraySlice_l173_252;
  wire                when_ArraySlice_l165_253;
  wire                when_ArraySlice_l166_253;
  reg        [6:0]    _zz_when_ArraySlice_l173_253;
  wire       [5:0]    _zz_when_ArraySlice_l112_253;
  wire                when_ArraySlice_l112_253;
  wire                when_ArraySlice_l113_253;
  wire                when_ArraySlice_l118_253;
  wire                when_ArraySlice_l173_253;
  wire                when_ArraySlice_l165_254;
  wire                when_ArraySlice_l166_254;
  reg        [6:0]    _zz_when_ArraySlice_l173_254;
  wire       [5:0]    _zz_when_ArraySlice_l112_254;
  wire                when_ArraySlice_l112_254;
  wire                when_ArraySlice_l113_254;
  wire                when_ArraySlice_l118_254;
  wire                when_ArraySlice_l173_254;
  wire                when_ArraySlice_l165_255;
  wire                when_ArraySlice_l166_255;
  reg        [6:0]    _zz_when_ArraySlice_l173_255;
  wire       [5:0]    _zz_when_ArraySlice_l112_255;
  wire                when_ArraySlice_l112_255;
  wire                when_ArraySlice_l113_255;
  wire                when_ArraySlice_l118_255;
  wire                when_ArraySlice_l173_255;
  wire                when_ArraySlice_l311_1;
  wire                outputStreamArrayData_1_fire_12;
  wire                when_ArraySlice_l315_1;
  wire                when_ArraySlice_l301_1;
  wire                outputStreamArrayData_1_fire_13;
  wire                when_ArraySlice_l322_1;
  wire                when_ArraySlice_l240_2;
  wire                when_ArraySlice_l241_2;
  wire       [5:0]    _zz_outputStreamArrayData_2_valid_1;
  wire                _zz_io_pop_ready_10;
  wire       [63:0]   _zz_13;
  wire                when_ArraySlice_l246_2;
  wire                outputStreamArrayData_2_fire_7;
  wire                when_ArraySlice_l247_2;
  wire                when_ArraySlice_l248_2;
  wire                when_ArraySlice_l251_2;
  wire                outputStreamArrayData_2_fire_8;
  wire                when_ArraySlice_l256_2;
  wire                when_ArraySlice_l257_2;
  reg        [6:0]    _zz_when_ArraySlice_l259_2;
  wire       [5:0]    _zz_when_ArraySlice_l94_30;
  wire                when_ArraySlice_l94_30;
  wire                when_ArraySlice_l95_30;
  wire                when_ArraySlice_l99_30;
  wire                when_ArraySlice_l259_2;
  reg                 debug_0_32 /* verilator public */ ;
  reg                 debug_1_32 /* verilator public */ ;
  reg                 debug_2_32 /* verilator public */ ;
  reg                 debug_3_32 /* verilator public */ ;
  reg                 debug_4_32 /* verilator public */ ;
  reg                 debug_5_32 /* verilator public */ ;
  reg                 debug_6_32 /* verilator public */ ;
  reg                 debug_7_32 /* verilator public */ ;
  wire                when_ArraySlice_l165_256;
  wire                when_ArraySlice_l166_256;
  reg        [6:0]    _zz_when_ArraySlice_l173_256;
  wire       [5:0]    _zz_when_ArraySlice_l112_256;
  wire                when_ArraySlice_l112_256;
  wire                when_ArraySlice_l113_256;
  wire                when_ArraySlice_l118_256;
  wire                when_ArraySlice_l173_256;
  wire                when_ArraySlice_l165_257;
  wire                when_ArraySlice_l166_257;
  reg        [6:0]    _zz_when_ArraySlice_l173_257;
  wire       [5:0]    _zz_when_ArraySlice_l112_257;
  wire                when_ArraySlice_l112_257;
  wire                when_ArraySlice_l113_257;
  wire                when_ArraySlice_l118_257;
  wire                when_ArraySlice_l173_257;
  wire                when_ArraySlice_l165_258;
  wire                when_ArraySlice_l166_258;
  reg        [6:0]    _zz_when_ArraySlice_l173_258;
  wire       [5:0]    _zz_when_ArraySlice_l112_258;
  wire                when_ArraySlice_l112_258;
  wire                when_ArraySlice_l113_258;
  wire                when_ArraySlice_l118_258;
  wire                when_ArraySlice_l173_258;
  wire                when_ArraySlice_l165_259;
  wire                when_ArraySlice_l166_259;
  reg        [6:0]    _zz_when_ArraySlice_l173_259;
  wire       [5:0]    _zz_when_ArraySlice_l112_259;
  wire                when_ArraySlice_l112_259;
  wire                when_ArraySlice_l113_259;
  wire                when_ArraySlice_l118_259;
  wire                when_ArraySlice_l173_259;
  wire                when_ArraySlice_l165_260;
  wire                when_ArraySlice_l166_260;
  reg        [6:0]    _zz_when_ArraySlice_l173_260;
  wire       [5:0]    _zz_when_ArraySlice_l112_260;
  wire                when_ArraySlice_l112_260;
  wire                when_ArraySlice_l113_260;
  wire                when_ArraySlice_l118_260;
  wire                when_ArraySlice_l173_260;
  wire                when_ArraySlice_l165_261;
  wire                when_ArraySlice_l166_261;
  reg        [6:0]    _zz_when_ArraySlice_l173_261;
  wire       [5:0]    _zz_when_ArraySlice_l112_261;
  wire                when_ArraySlice_l112_261;
  wire                when_ArraySlice_l113_261;
  wire                when_ArraySlice_l118_261;
  wire                when_ArraySlice_l173_261;
  wire                when_ArraySlice_l165_262;
  wire                when_ArraySlice_l166_262;
  reg        [6:0]    _zz_when_ArraySlice_l173_262;
  wire       [5:0]    _zz_when_ArraySlice_l112_262;
  wire                when_ArraySlice_l112_262;
  wire                when_ArraySlice_l113_262;
  wire                when_ArraySlice_l118_262;
  wire                when_ArraySlice_l173_262;
  wire                when_ArraySlice_l165_263;
  wire                when_ArraySlice_l166_263;
  reg        [6:0]    _zz_when_ArraySlice_l173_263;
  wire       [5:0]    _zz_when_ArraySlice_l112_263;
  wire                when_ArraySlice_l112_263;
  wire                when_ArraySlice_l113_263;
  wire                when_ArraySlice_l118_263;
  wire                when_ArraySlice_l173_263;
  wire                when_ArraySlice_l265_2;
  wire                when_ArraySlice_l268_2;
  wire                when_ArraySlice_l272_2;
  wire                when_ArraySlice_l276_2;
  wire                outputStreamArrayData_2_fire_9;
  wire                when_ArraySlice_l277_2;
  reg        [6:0]    _zz_when_ArraySlice_l279_2;
  wire       [5:0]    _zz_when_ArraySlice_l94_31;
  wire                when_ArraySlice_l94_31;
  wire                when_ArraySlice_l95_31;
  wire                when_ArraySlice_l99_31;
  wire                when_ArraySlice_l279_2;
  reg                 debug_0_33 /* verilator public */ ;
  reg                 debug_1_33 /* verilator public */ ;
  reg                 debug_2_33 /* verilator public */ ;
  reg                 debug_3_33 /* verilator public */ ;
  reg                 debug_4_33 /* verilator public */ ;
  reg                 debug_5_33 /* verilator public */ ;
  reg                 debug_6_33 /* verilator public */ ;
  reg                 debug_7_33 /* verilator public */ ;
  wire                when_ArraySlice_l165_264;
  wire                when_ArraySlice_l166_264;
  reg        [6:0]    _zz_when_ArraySlice_l173_264;
  wire       [5:0]    _zz_when_ArraySlice_l112_264;
  wire                when_ArraySlice_l112_264;
  wire                when_ArraySlice_l113_264;
  wire                when_ArraySlice_l118_264;
  wire                when_ArraySlice_l173_264;
  wire                when_ArraySlice_l165_265;
  wire                when_ArraySlice_l166_265;
  reg        [6:0]    _zz_when_ArraySlice_l173_265;
  wire       [5:0]    _zz_when_ArraySlice_l112_265;
  wire                when_ArraySlice_l112_265;
  wire                when_ArraySlice_l113_265;
  wire                when_ArraySlice_l118_265;
  wire                when_ArraySlice_l173_265;
  wire                when_ArraySlice_l165_266;
  wire                when_ArraySlice_l166_266;
  reg        [6:0]    _zz_when_ArraySlice_l173_266;
  wire       [5:0]    _zz_when_ArraySlice_l112_266;
  wire                when_ArraySlice_l112_266;
  wire                when_ArraySlice_l113_266;
  wire                when_ArraySlice_l118_266;
  wire                when_ArraySlice_l173_266;
  wire                when_ArraySlice_l165_267;
  wire                when_ArraySlice_l166_267;
  reg        [6:0]    _zz_when_ArraySlice_l173_267;
  wire       [5:0]    _zz_when_ArraySlice_l112_267;
  wire                when_ArraySlice_l112_267;
  wire                when_ArraySlice_l113_267;
  wire                when_ArraySlice_l118_267;
  wire                when_ArraySlice_l173_267;
  wire                when_ArraySlice_l165_268;
  wire                when_ArraySlice_l166_268;
  reg        [6:0]    _zz_when_ArraySlice_l173_268;
  wire       [5:0]    _zz_when_ArraySlice_l112_268;
  wire                when_ArraySlice_l112_268;
  wire                when_ArraySlice_l113_268;
  wire                when_ArraySlice_l118_268;
  wire                when_ArraySlice_l173_268;
  wire                when_ArraySlice_l165_269;
  wire                when_ArraySlice_l166_269;
  reg        [6:0]    _zz_when_ArraySlice_l173_269;
  wire       [5:0]    _zz_when_ArraySlice_l112_269;
  wire                when_ArraySlice_l112_269;
  wire                when_ArraySlice_l113_269;
  wire                when_ArraySlice_l118_269;
  wire                when_ArraySlice_l173_269;
  wire                when_ArraySlice_l165_270;
  wire                when_ArraySlice_l166_270;
  reg        [6:0]    _zz_when_ArraySlice_l173_270;
  wire       [5:0]    _zz_when_ArraySlice_l112_270;
  wire                when_ArraySlice_l112_270;
  wire                when_ArraySlice_l113_270;
  wire                when_ArraySlice_l118_270;
  wire                when_ArraySlice_l173_270;
  wire                when_ArraySlice_l165_271;
  wire                when_ArraySlice_l166_271;
  reg        [6:0]    _zz_when_ArraySlice_l173_271;
  wire       [5:0]    _zz_when_ArraySlice_l112_271;
  wire                when_ArraySlice_l112_271;
  wire                when_ArraySlice_l113_271;
  wire                when_ArraySlice_l118_271;
  wire                when_ArraySlice_l173_271;
  wire                when_ArraySlice_l285_2;
  wire                when_ArraySlice_l288_2;
  wire                outputStreamArrayData_2_fire_10;
  wire                when_ArraySlice_l292_2;
  wire                outputStreamArrayData_2_fire_11;
  wire                when_ArraySlice_l303_2;
  reg        [6:0]    _zz_when_ArraySlice_l304_2;
  wire       [5:0]    _zz_when_ArraySlice_l94_32;
  wire                when_ArraySlice_l94_32;
  wire                when_ArraySlice_l95_32;
  wire                when_ArraySlice_l99_32;
  wire                when_ArraySlice_l304_2;
  reg                 debug_0_34 /* verilator public */ ;
  reg                 debug_1_34 /* verilator public */ ;
  reg                 debug_2_34 /* verilator public */ ;
  reg                 debug_3_34 /* verilator public */ ;
  reg                 debug_4_34 /* verilator public */ ;
  reg                 debug_5_34 /* verilator public */ ;
  reg                 debug_6_34 /* verilator public */ ;
  reg                 debug_7_34 /* verilator public */ ;
  wire                when_ArraySlice_l165_272;
  wire                when_ArraySlice_l166_272;
  reg        [6:0]    _zz_when_ArraySlice_l173_272;
  wire       [5:0]    _zz_when_ArraySlice_l112_272;
  wire                when_ArraySlice_l112_272;
  wire                when_ArraySlice_l113_272;
  wire                when_ArraySlice_l118_272;
  wire                when_ArraySlice_l173_272;
  wire                when_ArraySlice_l165_273;
  wire                when_ArraySlice_l166_273;
  reg        [6:0]    _zz_when_ArraySlice_l173_273;
  wire       [5:0]    _zz_when_ArraySlice_l112_273;
  wire                when_ArraySlice_l112_273;
  wire                when_ArraySlice_l113_273;
  wire                when_ArraySlice_l118_273;
  wire                when_ArraySlice_l173_273;
  wire                when_ArraySlice_l165_274;
  wire                when_ArraySlice_l166_274;
  reg        [6:0]    _zz_when_ArraySlice_l173_274;
  wire       [5:0]    _zz_when_ArraySlice_l112_274;
  wire                when_ArraySlice_l112_274;
  wire                when_ArraySlice_l113_274;
  wire                when_ArraySlice_l118_274;
  wire                when_ArraySlice_l173_274;
  wire                when_ArraySlice_l165_275;
  wire                when_ArraySlice_l166_275;
  reg        [6:0]    _zz_when_ArraySlice_l173_275;
  wire       [5:0]    _zz_when_ArraySlice_l112_275;
  wire                when_ArraySlice_l112_275;
  wire                when_ArraySlice_l113_275;
  wire                when_ArraySlice_l118_275;
  wire                when_ArraySlice_l173_275;
  wire                when_ArraySlice_l165_276;
  wire                when_ArraySlice_l166_276;
  reg        [6:0]    _zz_when_ArraySlice_l173_276;
  wire       [5:0]    _zz_when_ArraySlice_l112_276;
  wire                when_ArraySlice_l112_276;
  wire                when_ArraySlice_l113_276;
  wire                when_ArraySlice_l118_276;
  wire                when_ArraySlice_l173_276;
  wire                when_ArraySlice_l165_277;
  wire                when_ArraySlice_l166_277;
  reg        [6:0]    _zz_when_ArraySlice_l173_277;
  wire       [5:0]    _zz_when_ArraySlice_l112_277;
  wire                when_ArraySlice_l112_277;
  wire                when_ArraySlice_l113_277;
  wire                when_ArraySlice_l118_277;
  wire                when_ArraySlice_l173_277;
  wire                when_ArraySlice_l165_278;
  wire                when_ArraySlice_l166_278;
  reg        [6:0]    _zz_when_ArraySlice_l173_278;
  wire       [5:0]    _zz_when_ArraySlice_l112_278;
  wire                when_ArraySlice_l112_278;
  wire                when_ArraySlice_l113_278;
  wire                when_ArraySlice_l118_278;
  wire                when_ArraySlice_l173_278;
  wire                when_ArraySlice_l165_279;
  wire                when_ArraySlice_l166_279;
  reg        [6:0]    _zz_when_ArraySlice_l173_279;
  wire       [5:0]    _zz_when_ArraySlice_l112_279;
  wire                when_ArraySlice_l112_279;
  wire                when_ArraySlice_l113_279;
  wire                when_ArraySlice_l118_279;
  wire                when_ArraySlice_l173_279;
  wire                when_ArraySlice_l311_2;
  wire                outputStreamArrayData_2_fire_12;
  wire                when_ArraySlice_l315_2;
  wire                when_ArraySlice_l301_2;
  wire                outputStreamArrayData_2_fire_13;
  wire                when_ArraySlice_l322_2;
  wire                when_ArraySlice_l240_3;
  wire                when_ArraySlice_l241_3;
  wire       [5:0]    _zz_outputStreamArrayData_3_valid_1;
  wire                _zz_io_pop_ready_11;
  wire       [63:0]   _zz_14;
  wire                when_ArraySlice_l246_3;
  wire                outputStreamArrayData_3_fire_7;
  wire                when_ArraySlice_l247_3;
  wire                when_ArraySlice_l248_3;
  wire                when_ArraySlice_l251_3;
  wire                outputStreamArrayData_3_fire_8;
  wire                when_ArraySlice_l256_3;
  wire                when_ArraySlice_l257_3;
  reg        [6:0]    _zz_when_ArraySlice_l259_3;
  wire       [5:0]    _zz_when_ArraySlice_l94_33;
  wire                when_ArraySlice_l94_33;
  wire                when_ArraySlice_l95_33;
  wire                when_ArraySlice_l99_33;
  wire                when_ArraySlice_l259_3;
  reg                 debug_0_35 /* verilator public */ ;
  reg                 debug_1_35 /* verilator public */ ;
  reg                 debug_2_35 /* verilator public */ ;
  reg                 debug_3_35 /* verilator public */ ;
  reg                 debug_4_35 /* verilator public */ ;
  reg                 debug_5_35 /* verilator public */ ;
  reg                 debug_6_35 /* verilator public */ ;
  reg                 debug_7_35 /* verilator public */ ;
  wire                when_ArraySlice_l165_280;
  wire                when_ArraySlice_l166_280;
  reg        [6:0]    _zz_when_ArraySlice_l173_280;
  wire       [5:0]    _zz_when_ArraySlice_l112_280;
  wire                when_ArraySlice_l112_280;
  wire                when_ArraySlice_l113_280;
  wire                when_ArraySlice_l118_280;
  wire                when_ArraySlice_l173_280;
  wire                when_ArraySlice_l165_281;
  wire                when_ArraySlice_l166_281;
  reg        [6:0]    _zz_when_ArraySlice_l173_281;
  wire       [5:0]    _zz_when_ArraySlice_l112_281;
  wire                when_ArraySlice_l112_281;
  wire                when_ArraySlice_l113_281;
  wire                when_ArraySlice_l118_281;
  wire                when_ArraySlice_l173_281;
  wire                when_ArraySlice_l165_282;
  wire                when_ArraySlice_l166_282;
  reg        [6:0]    _zz_when_ArraySlice_l173_282;
  wire       [5:0]    _zz_when_ArraySlice_l112_282;
  wire                when_ArraySlice_l112_282;
  wire                when_ArraySlice_l113_282;
  wire                when_ArraySlice_l118_282;
  wire                when_ArraySlice_l173_282;
  wire                when_ArraySlice_l165_283;
  wire                when_ArraySlice_l166_283;
  reg        [6:0]    _zz_when_ArraySlice_l173_283;
  wire       [5:0]    _zz_when_ArraySlice_l112_283;
  wire                when_ArraySlice_l112_283;
  wire                when_ArraySlice_l113_283;
  wire                when_ArraySlice_l118_283;
  wire                when_ArraySlice_l173_283;
  wire                when_ArraySlice_l165_284;
  wire                when_ArraySlice_l166_284;
  reg        [6:0]    _zz_when_ArraySlice_l173_284;
  wire       [5:0]    _zz_when_ArraySlice_l112_284;
  wire                when_ArraySlice_l112_284;
  wire                when_ArraySlice_l113_284;
  wire                when_ArraySlice_l118_284;
  wire                when_ArraySlice_l173_284;
  wire                when_ArraySlice_l165_285;
  wire                when_ArraySlice_l166_285;
  reg        [6:0]    _zz_when_ArraySlice_l173_285;
  wire       [5:0]    _zz_when_ArraySlice_l112_285;
  wire                when_ArraySlice_l112_285;
  wire                when_ArraySlice_l113_285;
  wire                when_ArraySlice_l118_285;
  wire                when_ArraySlice_l173_285;
  wire                when_ArraySlice_l165_286;
  wire                when_ArraySlice_l166_286;
  reg        [6:0]    _zz_when_ArraySlice_l173_286;
  wire       [5:0]    _zz_when_ArraySlice_l112_286;
  wire                when_ArraySlice_l112_286;
  wire                when_ArraySlice_l113_286;
  wire                when_ArraySlice_l118_286;
  wire                when_ArraySlice_l173_286;
  wire                when_ArraySlice_l165_287;
  wire                when_ArraySlice_l166_287;
  reg        [6:0]    _zz_when_ArraySlice_l173_287;
  wire       [5:0]    _zz_when_ArraySlice_l112_287;
  wire                when_ArraySlice_l112_287;
  wire                when_ArraySlice_l113_287;
  wire                when_ArraySlice_l118_287;
  wire                when_ArraySlice_l173_287;
  wire                when_ArraySlice_l265_3;
  wire                when_ArraySlice_l268_3;
  wire                when_ArraySlice_l272_3;
  wire                when_ArraySlice_l276_3;
  wire                outputStreamArrayData_3_fire_9;
  wire                when_ArraySlice_l277_3;
  reg        [6:0]    _zz_when_ArraySlice_l279_3;
  wire       [5:0]    _zz_when_ArraySlice_l94_34;
  wire                when_ArraySlice_l94_34;
  wire                when_ArraySlice_l95_34;
  wire                when_ArraySlice_l99_34;
  wire                when_ArraySlice_l279_3;
  reg                 debug_0_36 /* verilator public */ ;
  reg                 debug_1_36 /* verilator public */ ;
  reg                 debug_2_36 /* verilator public */ ;
  reg                 debug_3_36 /* verilator public */ ;
  reg                 debug_4_36 /* verilator public */ ;
  reg                 debug_5_36 /* verilator public */ ;
  reg                 debug_6_36 /* verilator public */ ;
  reg                 debug_7_36 /* verilator public */ ;
  wire                when_ArraySlice_l165_288;
  wire                when_ArraySlice_l166_288;
  reg        [6:0]    _zz_when_ArraySlice_l173_288;
  wire       [5:0]    _zz_when_ArraySlice_l112_288;
  wire                when_ArraySlice_l112_288;
  wire                when_ArraySlice_l113_288;
  wire                when_ArraySlice_l118_288;
  wire                when_ArraySlice_l173_288;
  wire                when_ArraySlice_l165_289;
  wire                when_ArraySlice_l166_289;
  reg        [6:0]    _zz_when_ArraySlice_l173_289;
  wire       [5:0]    _zz_when_ArraySlice_l112_289;
  wire                when_ArraySlice_l112_289;
  wire                when_ArraySlice_l113_289;
  wire                when_ArraySlice_l118_289;
  wire                when_ArraySlice_l173_289;
  wire                when_ArraySlice_l165_290;
  wire                when_ArraySlice_l166_290;
  reg        [6:0]    _zz_when_ArraySlice_l173_290;
  wire       [5:0]    _zz_when_ArraySlice_l112_290;
  wire                when_ArraySlice_l112_290;
  wire                when_ArraySlice_l113_290;
  wire                when_ArraySlice_l118_290;
  wire                when_ArraySlice_l173_290;
  wire                when_ArraySlice_l165_291;
  wire                when_ArraySlice_l166_291;
  reg        [6:0]    _zz_when_ArraySlice_l173_291;
  wire       [5:0]    _zz_when_ArraySlice_l112_291;
  wire                when_ArraySlice_l112_291;
  wire                when_ArraySlice_l113_291;
  wire                when_ArraySlice_l118_291;
  wire                when_ArraySlice_l173_291;
  wire                when_ArraySlice_l165_292;
  wire                when_ArraySlice_l166_292;
  reg        [6:0]    _zz_when_ArraySlice_l173_292;
  wire       [5:0]    _zz_when_ArraySlice_l112_292;
  wire                when_ArraySlice_l112_292;
  wire                when_ArraySlice_l113_292;
  wire                when_ArraySlice_l118_292;
  wire                when_ArraySlice_l173_292;
  wire                when_ArraySlice_l165_293;
  wire                when_ArraySlice_l166_293;
  reg        [6:0]    _zz_when_ArraySlice_l173_293;
  wire       [5:0]    _zz_when_ArraySlice_l112_293;
  wire                when_ArraySlice_l112_293;
  wire                when_ArraySlice_l113_293;
  wire                when_ArraySlice_l118_293;
  wire                when_ArraySlice_l173_293;
  wire                when_ArraySlice_l165_294;
  wire                when_ArraySlice_l166_294;
  reg        [6:0]    _zz_when_ArraySlice_l173_294;
  wire       [5:0]    _zz_when_ArraySlice_l112_294;
  wire                when_ArraySlice_l112_294;
  wire                when_ArraySlice_l113_294;
  wire                when_ArraySlice_l118_294;
  wire                when_ArraySlice_l173_294;
  wire                when_ArraySlice_l165_295;
  wire                when_ArraySlice_l166_295;
  reg        [6:0]    _zz_when_ArraySlice_l173_295;
  wire       [5:0]    _zz_when_ArraySlice_l112_295;
  wire                when_ArraySlice_l112_295;
  wire                when_ArraySlice_l113_295;
  wire                when_ArraySlice_l118_295;
  wire                when_ArraySlice_l173_295;
  wire                when_ArraySlice_l285_3;
  wire                when_ArraySlice_l288_3;
  wire                outputStreamArrayData_3_fire_10;
  wire                when_ArraySlice_l292_3;
  wire                outputStreamArrayData_3_fire_11;
  wire                when_ArraySlice_l303_3;
  reg        [6:0]    _zz_when_ArraySlice_l304_3;
  wire       [5:0]    _zz_when_ArraySlice_l94_35;
  wire                when_ArraySlice_l94_35;
  wire                when_ArraySlice_l95_35;
  wire                when_ArraySlice_l99_35;
  wire                when_ArraySlice_l304_3;
  reg                 debug_0_37 /* verilator public */ ;
  reg                 debug_1_37 /* verilator public */ ;
  reg                 debug_2_37 /* verilator public */ ;
  reg                 debug_3_37 /* verilator public */ ;
  reg                 debug_4_37 /* verilator public */ ;
  reg                 debug_5_37 /* verilator public */ ;
  reg                 debug_6_37 /* verilator public */ ;
  reg                 debug_7_37 /* verilator public */ ;
  wire                when_ArraySlice_l165_296;
  wire                when_ArraySlice_l166_296;
  reg        [6:0]    _zz_when_ArraySlice_l173_296;
  wire       [5:0]    _zz_when_ArraySlice_l112_296;
  wire                when_ArraySlice_l112_296;
  wire                when_ArraySlice_l113_296;
  wire                when_ArraySlice_l118_296;
  wire                when_ArraySlice_l173_296;
  wire                when_ArraySlice_l165_297;
  wire                when_ArraySlice_l166_297;
  reg        [6:0]    _zz_when_ArraySlice_l173_297;
  wire       [5:0]    _zz_when_ArraySlice_l112_297;
  wire                when_ArraySlice_l112_297;
  wire                when_ArraySlice_l113_297;
  wire                when_ArraySlice_l118_297;
  wire                when_ArraySlice_l173_297;
  wire                when_ArraySlice_l165_298;
  wire                when_ArraySlice_l166_298;
  reg        [6:0]    _zz_when_ArraySlice_l173_298;
  wire       [5:0]    _zz_when_ArraySlice_l112_298;
  wire                when_ArraySlice_l112_298;
  wire                when_ArraySlice_l113_298;
  wire                when_ArraySlice_l118_298;
  wire                when_ArraySlice_l173_298;
  wire                when_ArraySlice_l165_299;
  wire                when_ArraySlice_l166_299;
  reg        [6:0]    _zz_when_ArraySlice_l173_299;
  wire       [5:0]    _zz_when_ArraySlice_l112_299;
  wire                when_ArraySlice_l112_299;
  wire                when_ArraySlice_l113_299;
  wire                when_ArraySlice_l118_299;
  wire                when_ArraySlice_l173_299;
  wire                when_ArraySlice_l165_300;
  wire                when_ArraySlice_l166_300;
  reg        [6:0]    _zz_when_ArraySlice_l173_300;
  wire       [5:0]    _zz_when_ArraySlice_l112_300;
  wire                when_ArraySlice_l112_300;
  wire                when_ArraySlice_l113_300;
  wire                when_ArraySlice_l118_300;
  wire                when_ArraySlice_l173_300;
  wire                when_ArraySlice_l165_301;
  wire                when_ArraySlice_l166_301;
  reg        [6:0]    _zz_when_ArraySlice_l173_301;
  wire       [5:0]    _zz_when_ArraySlice_l112_301;
  wire                when_ArraySlice_l112_301;
  wire                when_ArraySlice_l113_301;
  wire                when_ArraySlice_l118_301;
  wire                when_ArraySlice_l173_301;
  wire                when_ArraySlice_l165_302;
  wire                when_ArraySlice_l166_302;
  reg        [6:0]    _zz_when_ArraySlice_l173_302;
  wire       [5:0]    _zz_when_ArraySlice_l112_302;
  wire                when_ArraySlice_l112_302;
  wire                when_ArraySlice_l113_302;
  wire                when_ArraySlice_l118_302;
  wire                when_ArraySlice_l173_302;
  wire                when_ArraySlice_l165_303;
  wire                when_ArraySlice_l166_303;
  reg        [6:0]    _zz_when_ArraySlice_l173_303;
  wire       [5:0]    _zz_when_ArraySlice_l112_303;
  wire                when_ArraySlice_l112_303;
  wire                when_ArraySlice_l113_303;
  wire                when_ArraySlice_l118_303;
  wire                when_ArraySlice_l173_303;
  wire                when_ArraySlice_l311_3;
  wire                outputStreamArrayData_3_fire_12;
  wire                when_ArraySlice_l315_3;
  wire                when_ArraySlice_l301_3;
  wire                outputStreamArrayData_3_fire_13;
  wire                when_ArraySlice_l322_3;
  wire                when_ArraySlice_l240_4;
  wire                when_ArraySlice_l241_4;
  wire       [5:0]    _zz_outputStreamArrayData_4_valid_1;
  wire                _zz_io_pop_ready_12;
  wire       [63:0]   _zz_15;
  wire                when_ArraySlice_l246_4;
  wire                outputStreamArrayData_4_fire_7;
  wire                when_ArraySlice_l247_4;
  wire                when_ArraySlice_l248_4;
  wire                when_ArraySlice_l251_4;
  wire                outputStreamArrayData_4_fire_8;
  wire                when_ArraySlice_l256_4;
  wire                when_ArraySlice_l257_4;
  reg        [6:0]    _zz_when_ArraySlice_l259_4;
  wire       [5:0]    _zz_when_ArraySlice_l94_36;
  wire                when_ArraySlice_l94_36;
  wire                when_ArraySlice_l95_36;
  wire                when_ArraySlice_l99_36;
  wire                when_ArraySlice_l259_4;
  reg                 debug_0_38 /* verilator public */ ;
  reg                 debug_1_38 /* verilator public */ ;
  reg                 debug_2_38 /* verilator public */ ;
  reg                 debug_3_38 /* verilator public */ ;
  reg                 debug_4_38 /* verilator public */ ;
  reg                 debug_5_38 /* verilator public */ ;
  reg                 debug_6_38 /* verilator public */ ;
  reg                 debug_7_38 /* verilator public */ ;
  wire                when_ArraySlice_l165_304;
  wire                when_ArraySlice_l166_304;
  reg        [6:0]    _zz_when_ArraySlice_l173_304;
  wire       [5:0]    _zz_when_ArraySlice_l112_304;
  wire                when_ArraySlice_l112_304;
  wire                when_ArraySlice_l113_304;
  wire                when_ArraySlice_l118_304;
  wire                when_ArraySlice_l173_304;
  wire                when_ArraySlice_l165_305;
  wire                when_ArraySlice_l166_305;
  reg        [6:0]    _zz_when_ArraySlice_l173_305;
  wire       [5:0]    _zz_when_ArraySlice_l112_305;
  wire                when_ArraySlice_l112_305;
  wire                when_ArraySlice_l113_305;
  wire                when_ArraySlice_l118_305;
  wire                when_ArraySlice_l173_305;
  wire                when_ArraySlice_l165_306;
  wire                when_ArraySlice_l166_306;
  reg        [6:0]    _zz_when_ArraySlice_l173_306;
  wire       [5:0]    _zz_when_ArraySlice_l112_306;
  wire                when_ArraySlice_l112_306;
  wire                when_ArraySlice_l113_306;
  wire                when_ArraySlice_l118_306;
  wire                when_ArraySlice_l173_306;
  wire                when_ArraySlice_l165_307;
  wire                when_ArraySlice_l166_307;
  reg        [6:0]    _zz_when_ArraySlice_l173_307;
  wire       [5:0]    _zz_when_ArraySlice_l112_307;
  wire                when_ArraySlice_l112_307;
  wire                when_ArraySlice_l113_307;
  wire                when_ArraySlice_l118_307;
  wire                when_ArraySlice_l173_307;
  wire                when_ArraySlice_l165_308;
  wire                when_ArraySlice_l166_308;
  reg        [6:0]    _zz_when_ArraySlice_l173_308;
  wire       [5:0]    _zz_when_ArraySlice_l112_308;
  wire                when_ArraySlice_l112_308;
  wire                when_ArraySlice_l113_308;
  wire                when_ArraySlice_l118_308;
  wire                when_ArraySlice_l173_308;
  wire                when_ArraySlice_l165_309;
  wire                when_ArraySlice_l166_309;
  reg        [6:0]    _zz_when_ArraySlice_l173_309;
  wire       [5:0]    _zz_when_ArraySlice_l112_309;
  wire                when_ArraySlice_l112_309;
  wire                when_ArraySlice_l113_309;
  wire                when_ArraySlice_l118_309;
  wire                when_ArraySlice_l173_309;
  wire                when_ArraySlice_l165_310;
  wire                when_ArraySlice_l166_310;
  reg        [6:0]    _zz_when_ArraySlice_l173_310;
  wire       [5:0]    _zz_when_ArraySlice_l112_310;
  wire                when_ArraySlice_l112_310;
  wire                when_ArraySlice_l113_310;
  wire                when_ArraySlice_l118_310;
  wire                when_ArraySlice_l173_310;
  wire                when_ArraySlice_l165_311;
  wire                when_ArraySlice_l166_311;
  reg        [6:0]    _zz_when_ArraySlice_l173_311;
  wire       [5:0]    _zz_when_ArraySlice_l112_311;
  wire                when_ArraySlice_l112_311;
  wire                when_ArraySlice_l113_311;
  wire                when_ArraySlice_l118_311;
  wire                when_ArraySlice_l173_311;
  wire                when_ArraySlice_l265_4;
  wire                when_ArraySlice_l268_4;
  wire                when_ArraySlice_l272_4;
  wire                when_ArraySlice_l276_4;
  wire                outputStreamArrayData_4_fire_9;
  wire                when_ArraySlice_l277_4;
  reg        [6:0]    _zz_when_ArraySlice_l279_4;
  wire       [5:0]    _zz_when_ArraySlice_l94_37;
  wire                when_ArraySlice_l94_37;
  wire                when_ArraySlice_l95_37;
  wire                when_ArraySlice_l99_37;
  wire                when_ArraySlice_l279_4;
  reg                 debug_0_39 /* verilator public */ ;
  reg                 debug_1_39 /* verilator public */ ;
  reg                 debug_2_39 /* verilator public */ ;
  reg                 debug_3_39 /* verilator public */ ;
  reg                 debug_4_39 /* verilator public */ ;
  reg                 debug_5_39 /* verilator public */ ;
  reg                 debug_6_39 /* verilator public */ ;
  reg                 debug_7_39 /* verilator public */ ;
  wire                when_ArraySlice_l165_312;
  wire                when_ArraySlice_l166_312;
  reg        [6:0]    _zz_when_ArraySlice_l173_312;
  wire       [5:0]    _zz_when_ArraySlice_l112_312;
  wire                when_ArraySlice_l112_312;
  wire                when_ArraySlice_l113_312;
  wire                when_ArraySlice_l118_312;
  wire                when_ArraySlice_l173_312;
  wire                when_ArraySlice_l165_313;
  wire                when_ArraySlice_l166_313;
  reg        [6:0]    _zz_when_ArraySlice_l173_313;
  wire       [5:0]    _zz_when_ArraySlice_l112_313;
  wire                when_ArraySlice_l112_313;
  wire                when_ArraySlice_l113_313;
  wire                when_ArraySlice_l118_313;
  wire                when_ArraySlice_l173_313;
  wire                when_ArraySlice_l165_314;
  wire                when_ArraySlice_l166_314;
  reg        [6:0]    _zz_when_ArraySlice_l173_314;
  wire       [5:0]    _zz_when_ArraySlice_l112_314;
  wire                when_ArraySlice_l112_314;
  wire                when_ArraySlice_l113_314;
  wire                when_ArraySlice_l118_314;
  wire                when_ArraySlice_l173_314;
  wire                when_ArraySlice_l165_315;
  wire                when_ArraySlice_l166_315;
  reg        [6:0]    _zz_when_ArraySlice_l173_315;
  wire       [5:0]    _zz_when_ArraySlice_l112_315;
  wire                when_ArraySlice_l112_315;
  wire                when_ArraySlice_l113_315;
  wire                when_ArraySlice_l118_315;
  wire                when_ArraySlice_l173_315;
  wire                when_ArraySlice_l165_316;
  wire                when_ArraySlice_l166_316;
  reg        [6:0]    _zz_when_ArraySlice_l173_316;
  wire       [5:0]    _zz_when_ArraySlice_l112_316;
  wire                when_ArraySlice_l112_316;
  wire                when_ArraySlice_l113_316;
  wire                when_ArraySlice_l118_316;
  wire                when_ArraySlice_l173_316;
  wire                when_ArraySlice_l165_317;
  wire                when_ArraySlice_l166_317;
  reg        [6:0]    _zz_when_ArraySlice_l173_317;
  wire       [5:0]    _zz_when_ArraySlice_l112_317;
  wire                when_ArraySlice_l112_317;
  wire                when_ArraySlice_l113_317;
  wire                when_ArraySlice_l118_317;
  wire                when_ArraySlice_l173_317;
  wire                when_ArraySlice_l165_318;
  wire                when_ArraySlice_l166_318;
  reg        [6:0]    _zz_when_ArraySlice_l173_318;
  wire       [5:0]    _zz_when_ArraySlice_l112_318;
  wire                when_ArraySlice_l112_318;
  wire                when_ArraySlice_l113_318;
  wire                when_ArraySlice_l118_318;
  wire                when_ArraySlice_l173_318;
  wire                when_ArraySlice_l165_319;
  wire                when_ArraySlice_l166_319;
  reg        [6:0]    _zz_when_ArraySlice_l173_319;
  wire       [5:0]    _zz_when_ArraySlice_l112_319;
  wire                when_ArraySlice_l112_319;
  wire                when_ArraySlice_l113_319;
  wire                when_ArraySlice_l118_319;
  wire                when_ArraySlice_l173_319;
  wire                when_ArraySlice_l285_4;
  wire                when_ArraySlice_l288_4;
  wire                outputStreamArrayData_4_fire_10;
  wire                when_ArraySlice_l292_4;
  wire                outputStreamArrayData_4_fire_11;
  wire                when_ArraySlice_l303_4;
  reg        [6:0]    _zz_when_ArraySlice_l304_4;
  wire       [5:0]    _zz_when_ArraySlice_l94_38;
  wire                when_ArraySlice_l94_38;
  wire                when_ArraySlice_l95_38;
  wire                when_ArraySlice_l99_38;
  wire                when_ArraySlice_l304_4;
  reg                 debug_0_40 /* verilator public */ ;
  reg                 debug_1_40 /* verilator public */ ;
  reg                 debug_2_40 /* verilator public */ ;
  reg                 debug_3_40 /* verilator public */ ;
  reg                 debug_4_40 /* verilator public */ ;
  reg                 debug_5_40 /* verilator public */ ;
  reg                 debug_6_40 /* verilator public */ ;
  reg                 debug_7_40 /* verilator public */ ;
  wire                when_ArraySlice_l165_320;
  wire                when_ArraySlice_l166_320;
  reg        [6:0]    _zz_when_ArraySlice_l173_320;
  wire       [5:0]    _zz_when_ArraySlice_l112_320;
  wire                when_ArraySlice_l112_320;
  wire                when_ArraySlice_l113_320;
  wire                when_ArraySlice_l118_320;
  wire                when_ArraySlice_l173_320;
  wire                when_ArraySlice_l165_321;
  wire                when_ArraySlice_l166_321;
  reg        [6:0]    _zz_when_ArraySlice_l173_321;
  wire       [5:0]    _zz_when_ArraySlice_l112_321;
  wire                when_ArraySlice_l112_321;
  wire                when_ArraySlice_l113_321;
  wire                when_ArraySlice_l118_321;
  wire                when_ArraySlice_l173_321;
  wire                when_ArraySlice_l165_322;
  wire                when_ArraySlice_l166_322;
  reg        [6:0]    _zz_when_ArraySlice_l173_322;
  wire       [5:0]    _zz_when_ArraySlice_l112_322;
  wire                when_ArraySlice_l112_322;
  wire                when_ArraySlice_l113_322;
  wire                when_ArraySlice_l118_322;
  wire                when_ArraySlice_l173_322;
  wire                when_ArraySlice_l165_323;
  wire                when_ArraySlice_l166_323;
  reg        [6:0]    _zz_when_ArraySlice_l173_323;
  wire       [5:0]    _zz_when_ArraySlice_l112_323;
  wire                when_ArraySlice_l112_323;
  wire                when_ArraySlice_l113_323;
  wire                when_ArraySlice_l118_323;
  wire                when_ArraySlice_l173_323;
  wire                when_ArraySlice_l165_324;
  wire                when_ArraySlice_l166_324;
  reg        [6:0]    _zz_when_ArraySlice_l173_324;
  wire       [5:0]    _zz_when_ArraySlice_l112_324;
  wire                when_ArraySlice_l112_324;
  wire                when_ArraySlice_l113_324;
  wire                when_ArraySlice_l118_324;
  wire                when_ArraySlice_l173_324;
  wire                when_ArraySlice_l165_325;
  wire                when_ArraySlice_l166_325;
  reg        [6:0]    _zz_when_ArraySlice_l173_325;
  wire       [5:0]    _zz_when_ArraySlice_l112_325;
  wire                when_ArraySlice_l112_325;
  wire                when_ArraySlice_l113_325;
  wire                when_ArraySlice_l118_325;
  wire                when_ArraySlice_l173_325;
  wire                when_ArraySlice_l165_326;
  wire                when_ArraySlice_l166_326;
  reg        [6:0]    _zz_when_ArraySlice_l173_326;
  wire       [5:0]    _zz_when_ArraySlice_l112_326;
  wire                when_ArraySlice_l112_326;
  wire                when_ArraySlice_l113_326;
  wire                when_ArraySlice_l118_326;
  wire                when_ArraySlice_l173_326;
  wire                when_ArraySlice_l165_327;
  wire                when_ArraySlice_l166_327;
  reg        [6:0]    _zz_when_ArraySlice_l173_327;
  wire       [5:0]    _zz_when_ArraySlice_l112_327;
  wire                when_ArraySlice_l112_327;
  wire                when_ArraySlice_l113_327;
  wire                when_ArraySlice_l118_327;
  wire                when_ArraySlice_l173_327;
  wire                when_ArraySlice_l311_4;
  wire                outputStreamArrayData_4_fire_12;
  wire                when_ArraySlice_l315_4;
  wire                when_ArraySlice_l301_4;
  wire                outputStreamArrayData_4_fire_13;
  wire                when_ArraySlice_l322_4;
  wire                when_ArraySlice_l240_5;
  wire                when_ArraySlice_l241_5;
  wire       [5:0]    _zz_outputStreamArrayData_5_valid_1;
  wire                _zz_io_pop_ready_13;
  wire       [63:0]   _zz_16;
  wire                when_ArraySlice_l246_5;
  wire                outputStreamArrayData_5_fire_7;
  wire                when_ArraySlice_l247_5;
  wire                when_ArraySlice_l248_5;
  wire                when_ArraySlice_l251_5;
  wire                outputStreamArrayData_5_fire_8;
  wire                when_ArraySlice_l256_5;
  wire                when_ArraySlice_l257_5;
  reg        [6:0]    _zz_when_ArraySlice_l259_5;
  wire       [5:0]    _zz_when_ArraySlice_l94_39;
  wire                when_ArraySlice_l94_39;
  wire                when_ArraySlice_l95_39;
  wire                when_ArraySlice_l99_39;
  wire                when_ArraySlice_l259_5;
  reg                 debug_0_41 /* verilator public */ ;
  reg                 debug_1_41 /* verilator public */ ;
  reg                 debug_2_41 /* verilator public */ ;
  reg                 debug_3_41 /* verilator public */ ;
  reg                 debug_4_41 /* verilator public */ ;
  reg                 debug_5_41 /* verilator public */ ;
  reg                 debug_6_41 /* verilator public */ ;
  reg                 debug_7_41 /* verilator public */ ;
  wire                when_ArraySlice_l165_328;
  wire                when_ArraySlice_l166_328;
  reg        [6:0]    _zz_when_ArraySlice_l173_328;
  wire       [5:0]    _zz_when_ArraySlice_l112_328;
  wire                when_ArraySlice_l112_328;
  wire                when_ArraySlice_l113_328;
  wire                when_ArraySlice_l118_328;
  wire                when_ArraySlice_l173_328;
  wire                when_ArraySlice_l165_329;
  wire                when_ArraySlice_l166_329;
  reg        [6:0]    _zz_when_ArraySlice_l173_329;
  wire       [5:0]    _zz_when_ArraySlice_l112_329;
  wire                when_ArraySlice_l112_329;
  wire                when_ArraySlice_l113_329;
  wire                when_ArraySlice_l118_329;
  wire                when_ArraySlice_l173_329;
  wire                when_ArraySlice_l165_330;
  wire                when_ArraySlice_l166_330;
  reg        [6:0]    _zz_when_ArraySlice_l173_330;
  wire       [5:0]    _zz_when_ArraySlice_l112_330;
  wire                when_ArraySlice_l112_330;
  wire                when_ArraySlice_l113_330;
  wire                when_ArraySlice_l118_330;
  wire                when_ArraySlice_l173_330;
  wire                when_ArraySlice_l165_331;
  wire                when_ArraySlice_l166_331;
  reg        [6:0]    _zz_when_ArraySlice_l173_331;
  wire       [5:0]    _zz_when_ArraySlice_l112_331;
  wire                when_ArraySlice_l112_331;
  wire                when_ArraySlice_l113_331;
  wire                when_ArraySlice_l118_331;
  wire                when_ArraySlice_l173_331;
  wire                when_ArraySlice_l165_332;
  wire                when_ArraySlice_l166_332;
  reg        [6:0]    _zz_when_ArraySlice_l173_332;
  wire       [5:0]    _zz_when_ArraySlice_l112_332;
  wire                when_ArraySlice_l112_332;
  wire                when_ArraySlice_l113_332;
  wire                when_ArraySlice_l118_332;
  wire                when_ArraySlice_l173_332;
  wire                when_ArraySlice_l165_333;
  wire                when_ArraySlice_l166_333;
  reg        [6:0]    _zz_when_ArraySlice_l173_333;
  wire       [5:0]    _zz_when_ArraySlice_l112_333;
  wire                when_ArraySlice_l112_333;
  wire                when_ArraySlice_l113_333;
  wire                when_ArraySlice_l118_333;
  wire                when_ArraySlice_l173_333;
  wire                when_ArraySlice_l165_334;
  wire                when_ArraySlice_l166_334;
  reg        [6:0]    _zz_when_ArraySlice_l173_334;
  wire       [5:0]    _zz_when_ArraySlice_l112_334;
  wire                when_ArraySlice_l112_334;
  wire                when_ArraySlice_l113_334;
  wire                when_ArraySlice_l118_334;
  wire                when_ArraySlice_l173_334;
  wire                when_ArraySlice_l165_335;
  wire                when_ArraySlice_l166_335;
  reg        [6:0]    _zz_when_ArraySlice_l173_335;
  wire       [5:0]    _zz_when_ArraySlice_l112_335;
  wire                when_ArraySlice_l112_335;
  wire                when_ArraySlice_l113_335;
  wire                when_ArraySlice_l118_335;
  wire                when_ArraySlice_l173_335;
  wire                when_ArraySlice_l265_5;
  wire                when_ArraySlice_l268_5;
  wire                when_ArraySlice_l272_5;
  wire                when_ArraySlice_l276_5;
  wire                outputStreamArrayData_5_fire_9;
  wire                when_ArraySlice_l277_5;
  reg        [6:0]    _zz_when_ArraySlice_l279_5;
  wire       [5:0]    _zz_when_ArraySlice_l94_40;
  wire                when_ArraySlice_l94_40;
  wire                when_ArraySlice_l95_40;
  wire                when_ArraySlice_l99_40;
  wire                when_ArraySlice_l279_5;
  reg                 debug_0_42 /* verilator public */ ;
  reg                 debug_1_42 /* verilator public */ ;
  reg                 debug_2_42 /* verilator public */ ;
  reg                 debug_3_42 /* verilator public */ ;
  reg                 debug_4_42 /* verilator public */ ;
  reg                 debug_5_42 /* verilator public */ ;
  reg                 debug_6_42 /* verilator public */ ;
  reg                 debug_7_42 /* verilator public */ ;
  wire                when_ArraySlice_l165_336;
  wire                when_ArraySlice_l166_336;
  reg        [6:0]    _zz_when_ArraySlice_l173_336;
  wire       [5:0]    _zz_when_ArraySlice_l112_336;
  wire                when_ArraySlice_l112_336;
  wire                when_ArraySlice_l113_336;
  wire                when_ArraySlice_l118_336;
  wire                when_ArraySlice_l173_336;
  wire                when_ArraySlice_l165_337;
  wire                when_ArraySlice_l166_337;
  reg        [6:0]    _zz_when_ArraySlice_l173_337;
  wire       [5:0]    _zz_when_ArraySlice_l112_337;
  wire                when_ArraySlice_l112_337;
  wire                when_ArraySlice_l113_337;
  wire                when_ArraySlice_l118_337;
  wire                when_ArraySlice_l173_337;
  wire                when_ArraySlice_l165_338;
  wire                when_ArraySlice_l166_338;
  reg        [6:0]    _zz_when_ArraySlice_l173_338;
  wire       [5:0]    _zz_when_ArraySlice_l112_338;
  wire                when_ArraySlice_l112_338;
  wire                when_ArraySlice_l113_338;
  wire                when_ArraySlice_l118_338;
  wire                when_ArraySlice_l173_338;
  wire                when_ArraySlice_l165_339;
  wire                when_ArraySlice_l166_339;
  reg        [6:0]    _zz_when_ArraySlice_l173_339;
  wire       [5:0]    _zz_when_ArraySlice_l112_339;
  wire                when_ArraySlice_l112_339;
  wire                when_ArraySlice_l113_339;
  wire                when_ArraySlice_l118_339;
  wire                when_ArraySlice_l173_339;
  wire                when_ArraySlice_l165_340;
  wire                when_ArraySlice_l166_340;
  reg        [6:0]    _zz_when_ArraySlice_l173_340;
  wire       [5:0]    _zz_when_ArraySlice_l112_340;
  wire                when_ArraySlice_l112_340;
  wire                when_ArraySlice_l113_340;
  wire                when_ArraySlice_l118_340;
  wire                when_ArraySlice_l173_340;
  wire                when_ArraySlice_l165_341;
  wire                when_ArraySlice_l166_341;
  reg        [6:0]    _zz_when_ArraySlice_l173_341;
  wire       [5:0]    _zz_when_ArraySlice_l112_341;
  wire                when_ArraySlice_l112_341;
  wire                when_ArraySlice_l113_341;
  wire                when_ArraySlice_l118_341;
  wire                when_ArraySlice_l173_341;
  wire                when_ArraySlice_l165_342;
  wire                when_ArraySlice_l166_342;
  reg        [6:0]    _zz_when_ArraySlice_l173_342;
  wire       [5:0]    _zz_when_ArraySlice_l112_342;
  wire                when_ArraySlice_l112_342;
  wire                when_ArraySlice_l113_342;
  wire                when_ArraySlice_l118_342;
  wire                when_ArraySlice_l173_342;
  wire                when_ArraySlice_l165_343;
  wire                when_ArraySlice_l166_343;
  reg        [6:0]    _zz_when_ArraySlice_l173_343;
  wire       [5:0]    _zz_when_ArraySlice_l112_343;
  wire                when_ArraySlice_l112_343;
  wire                when_ArraySlice_l113_343;
  wire                when_ArraySlice_l118_343;
  wire                when_ArraySlice_l173_343;
  wire                when_ArraySlice_l285_5;
  wire                when_ArraySlice_l288_5;
  wire                outputStreamArrayData_5_fire_10;
  wire                when_ArraySlice_l292_5;
  wire                outputStreamArrayData_5_fire_11;
  wire                when_ArraySlice_l303_5;
  reg        [6:0]    _zz_when_ArraySlice_l304_5;
  wire       [5:0]    _zz_when_ArraySlice_l94_41;
  wire                when_ArraySlice_l94_41;
  wire                when_ArraySlice_l95_41;
  wire                when_ArraySlice_l99_41;
  wire                when_ArraySlice_l304_5;
  reg                 debug_0_43 /* verilator public */ ;
  reg                 debug_1_43 /* verilator public */ ;
  reg                 debug_2_43 /* verilator public */ ;
  reg                 debug_3_43 /* verilator public */ ;
  reg                 debug_4_43 /* verilator public */ ;
  reg                 debug_5_43 /* verilator public */ ;
  reg                 debug_6_43 /* verilator public */ ;
  reg                 debug_7_43 /* verilator public */ ;
  wire                when_ArraySlice_l165_344;
  wire                when_ArraySlice_l166_344;
  reg        [6:0]    _zz_when_ArraySlice_l173_344;
  wire       [5:0]    _zz_when_ArraySlice_l112_344;
  wire                when_ArraySlice_l112_344;
  wire                when_ArraySlice_l113_344;
  wire                when_ArraySlice_l118_344;
  wire                when_ArraySlice_l173_344;
  wire                when_ArraySlice_l165_345;
  wire                when_ArraySlice_l166_345;
  reg        [6:0]    _zz_when_ArraySlice_l173_345;
  wire       [5:0]    _zz_when_ArraySlice_l112_345;
  wire                when_ArraySlice_l112_345;
  wire                when_ArraySlice_l113_345;
  wire                when_ArraySlice_l118_345;
  wire                when_ArraySlice_l173_345;
  wire                when_ArraySlice_l165_346;
  wire                when_ArraySlice_l166_346;
  reg        [6:0]    _zz_when_ArraySlice_l173_346;
  wire       [5:0]    _zz_when_ArraySlice_l112_346;
  wire                when_ArraySlice_l112_346;
  wire                when_ArraySlice_l113_346;
  wire                when_ArraySlice_l118_346;
  wire                when_ArraySlice_l173_346;
  wire                when_ArraySlice_l165_347;
  wire                when_ArraySlice_l166_347;
  reg        [6:0]    _zz_when_ArraySlice_l173_347;
  wire       [5:0]    _zz_when_ArraySlice_l112_347;
  wire                when_ArraySlice_l112_347;
  wire                when_ArraySlice_l113_347;
  wire                when_ArraySlice_l118_347;
  wire                when_ArraySlice_l173_347;
  wire                when_ArraySlice_l165_348;
  wire                when_ArraySlice_l166_348;
  reg        [6:0]    _zz_when_ArraySlice_l173_348;
  wire       [5:0]    _zz_when_ArraySlice_l112_348;
  wire                when_ArraySlice_l112_348;
  wire                when_ArraySlice_l113_348;
  wire                when_ArraySlice_l118_348;
  wire                when_ArraySlice_l173_348;
  wire                when_ArraySlice_l165_349;
  wire                when_ArraySlice_l166_349;
  reg        [6:0]    _zz_when_ArraySlice_l173_349;
  wire       [5:0]    _zz_when_ArraySlice_l112_349;
  wire                when_ArraySlice_l112_349;
  wire                when_ArraySlice_l113_349;
  wire                when_ArraySlice_l118_349;
  wire                when_ArraySlice_l173_349;
  wire                when_ArraySlice_l165_350;
  wire                when_ArraySlice_l166_350;
  reg        [6:0]    _zz_when_ArraySlice_l173_350;
  wire       [5:0]    _zz_when_ArraySlice_l112_350;
  wire                when_ArraySlice_l112_350;
  wire                when_ArraySlice_l113_350;
  wire                when_ArraySlice_l118_350;
  wire                when_ArraySlice_l173_350;
  wire                when_ArraySlice_l165_351;
  wire                when_ArraySlice_l166_351;
  reg        [6:0]    _zz_when_ArraySlice_l173_351;
  wire       [5:0]    _zz_when_ArraySlice_l112_351;
  wire                when_ArraySlice_l112_351;
  wire                when_ArraySlice_l113_351;
  wire                when_ArraySlice_l118_351;
  wire                when_ArraySlice_l173_351;
  wire                when_ArraySlice_l311_5;
  wire                outputStreamArrayData_5_fire_12;
  wire                when_ArraySlice_l315_5;
  wire                when_ArraySlice_l301_5;
  wire                outputStreamArrayData_5_fire_13;
  wire                when_ArraySlice_l322_5;
  wire                when_ArraySlice_l240_6;
  wire                when_ArraySlice_l241_6;
  wire       [5:0]    _zz_outputStreamArrayData_6_valid_1;
  wire                _zz_io_pop_ready_14;
  wire       [63:0]   _zz_17;
  wire                when_ArraySlice_l246_6;
  wire                outputStreamArrayData_6_fire_7;
  wire                when_ArraySlice_l247_6;
  wire                when_ArraySlice_l248_6;
  wire                when_ArraySlice_l251_6;
  wire                outputStreamArrayData_6_fire_8;
  wire                when_ArraySlice_l256_6;
  wire                when_ArraySlice_l257_6;
  reg        [6:0]    _zz_when_ArraySlice_l259_6;
  wire       [5:0]    _zz_when_ArraySlice_l94_42;
  wire                when_ArraySlice_l94_42;
  wire                when_ArraySlice_l95_42;
  wire                when_ArraySlice_l99_42;
  wire                when_ArraySlice_l259_6;
  reg                 debug_0_44 /* verilator public */ ;
  reg                 debug_1_44 /* verilator public */ ;
  reg                 debug_2_44 /* verilator public */ ;
  reg                 debug_3_44 /* verilator public */ ;
  reg                 debug_4_44 /* verilator public */ ;
  reg                 debug_5_44 /* verilator public */ ;
  reg                 debug_6_44 /* verilator public */ ;
  reg                 debug_7_44 /* verilator public */ ;
  wire                when_ArraySlice_l165_352;
  wire                when_ArraySlice_l166_352;
  reg        [6:0]    _zz_when_ArraySlice_l173_352;
  wire       [5:0]    _zz_when_ArraySlice_l112_352;
  wire                when_ArraySlice_l112_352;
  wire                when_ArraySlice_l113_352;
  wire                when_ArraySlice_l118_352;
  wire                when_ArraySlice_l173_352;
  wire                when_ArraySlice_l165_353;
  wire                when_ArraySlice_l166_353;
  reg        [6:0]    _zz_when_ArraySlice_l173_353;
  wire       [5:0]    _zz_when_ArraySlice_l112_353;
  wire                when_ArraySlice_l112_353;
  wire                when_ArraySlice_l113_353;
  wire                when_ArraySlice_l118_353;
  wire                when_ArraySlice_l173_353;
  wire                when_ArraySlice_l165_354;
  wire                when_ArraySlice_l166_354;
  reg        [6:0]    _zz_when_ArraySlice_l173_354;
  wire       [5:0]    _zz_when_ArraySlice_l112_354;
  wire                when_ArraySlice_l112_354;
  wire                when_ArraySlice_l113_354;
  wire                when_ArraySlice_l118_354;
  wire                when_ArraySlice_l173_354;
  wire                when_ArraySlice_l165_355;
  wire                when_ArraySlice_l166_355;
  reg        [6:0]    _zz_when_ArraySlice_l173_355;
  wire       [5:0]    _zz_when_ArraySlice_l112_355;
  wire                when_ArraySlice_l112_355;
  wire                when_ArraySlice_l113_355;
  wire                when_ArraySlice_l118_355;
  wire                when_ArraySlice_l173_355;
  wire                when_ArraySlice_l165_356;
  wire                when_ArraySlice_l166_356;
  reg        [6:0]    _zz_when_ArraySlice_l173_356;
  wire       [5:0]    _zz_when_ArraySlice_l112_356;
  wire                when_ArraySlice_l112_356;
  wire                when_ArraySlice_l113_356;
  wire                when_ArraySlice_l118_356;
  wire                when_ArraySlice_l173_356;
  wire                when_ArraySlice_l165_357;
  wire                when_ArraySlice_l166_357;
  reg        [6:0]    _zz_when_ArraySlice_l173_357;
  wire       [5:0]    _zz_when_ArraySlice_l112_357;
  wire                when_ArraySlice_l112_357;
  wire                when_ArraySlice_l113_357;
  wire                when_ArraySlice_l118_357;
  wire                when_ArraySlice_l173_357;
  wire                when_ArraySlice_l165_358;
  wire                when_ArraySlice_l166_358;
  reg        [6:0]    _zz_when_ArraySlice_l173_358;
  wire       [5:0]    _zz_when_ArraySlice_l112_358;
  wire                when_ArraySlice_l112_358;
  wire                when_ArraySlice_l113_358;
  wire                when_ArraySlice_l118_358;
  wire                when_ArraySlice_l173_358;
  wire                when_ArraySlice_l165_359;
  wire                when_ArraySlice_l166_359;
  reg        [6:0]    _zz_when_ArraySlice_l173_359;
  wire       [5:0]    _zz_when_ArraySlice_l112_359;
  wire                when_ArraySlice_l112_359;
  wire                when_ArraySlice_l113_359;
  wire                when_ArraySlice_l118_359;
  wire                when_ArraySlice_l173_359;
  wire                when_ArraySlice_l265_6;
  wire                when_ArraySlice_l268_6;
  wire                when_ArraySlice_l272_6;
  wire                when_ArraySlice_l276_6;
  wire                outputStreamArrayData_6_fire_9;
  wire                when_ArraySlice_l277_6;
  reg        [6:0]    _zz_when_ArraySlice_l279_6;
  wire       [5:0]    _zz_when_ArraySlice_l94_43;
  wire                when_ArraySlice_l94_43;
  wire                when_ArraySlice_l95_43;
  wire                when_ArraySlice_l99_43;
  wire                when_ArraySlice_l279_6;
  reg                 debug_0_45 /* verilator public */ ;
  reg                 debug_1_45 /* verilator public */ ;
  reg                 debug_2_45 /* verilator public */ ;
  reg                 debug_3_45 /* verilator public */ ;
  reg                 debug_4_45 /* verilator public */ ;
  reg                 debug_5_45 /* verilator public */ ;
  reg                 debug_6_45 /* verilator public */ ;
  reg                 debug_7_45 /* verilator public */ ;
  wire                when_ArraySlice_l165_360;
  wire                when_ArraySlice_l166_360;
  reg        [6:0]    _zz_when_ArraySlice_l173_360;
  wire       [5:0]    _zz_when_ArraySlice_l112_360;
  wire                when_ArraySlice_l112_360;
  wire                when_ArraySlice_l113_360;
  wire                when_ArraySlice_l118_360;
  wire                when_ArraySlice_l173_360;
  wire                when_ArraySlice_l165_361;
  wire                when_ArraySlice_l166_361;
  reg        [6:0]    _zz_when_ArraySlice_l173_361;
  wire       [5:0]    _zz_when_ArraySlice_l112_361;
  wire                when_ArraySlice_l112_361;
  wire                when_ArraySlice_l113_361;
  wire                when_ArraySlice_l118_361;
  wire                when_ArraySlice_l173_361;
  wire                when_ArraySlice_l165_362;
  wire                when_ArraySlice_l166_362;
  reg        [6:0]    _zz_when_ArraySlice_l173_362;
  wire       [5:0]    _zz_when_ArraySlice_l112_362;
  wire                when_ArraySlice_l112_362;
  wire                when_ArraySlice_l113_362;
  wire                when_ArraySlice_l118_362;
  wire                when_ArraySlice_l173_362;
  wire                when_ArraySlice_l165_363;
  wire                when_ArraySlice_l166_363;
  reg        [6:0]    _zz_when_ArraySlice_l173_363;
  wire       [5:0]    _zz_when_ArraySlice_l112_363;
  wire                when_ArraySlice_l112_363;
  wire                when_ArraySlice_l113_363;
  wire                when_ArraySlice_l118_363;
  wire                when_ArraySlice_l173_363;
  wire                when_ArraySlice_l165_364;
  wire                when_ArraySlice_l166_364;
  reg        [6:0]    _zz_when_ArraySlice_l173_364;
  wire       [5:0]    _zz_when_ArraySlice_l112_364;
  wire                when_ArraySlice_l112_364;
  wire                when_ArraySlice_l113_364;
  wire                when_ArraySlice_l118_364;
  wire                when_ArraySlice_l173_364;
  wire                when_ArraySlice_l165_365;
  wire                when_ArraySlice_l166_365;
  reg        [6:0]    _zz_when_ArraySlice_l173_365;
  wire       [5:0]    _zz_when_ArraySlice_l112_365;
  wire                when_ArraySlice_l112_365;
  wire                when_ArraySlice_l113_365;
  wire                when_ArraySlice_l118_365;
  wire                when_ArraySlice_l173_365;
  wire                when_ArraySlice_l165_366;
  wire                when_ArraySlice_l166_366;
  reg        [6:0]    _zz_when_ArraySlice_l173_366;
  wire       [5:0]    _zz_when_ArraySlice_l112_366;
  wire                when_ArraySlice_l112_366;
  wire                when_ArraySlice_l113_366;
  wire                when_ArraySlice_l118_366;
  wire                when_ArraySlice_l173_366;
  wire                when_ArraySlice_l165_367;
  wire                when_ArraySlice_l166_367;
  reg        [6:0]    _zz_when_ArraySlice_l173_367;
  wire       [5:0]    _zz_when_ArraySlice_l112_367;
  wire                when_ArraySlice_l112_367;
  wire                when_ArraySlice_l113_367;
  wire                when_ArraySlice_l118_367;
  wire                when_ArraySlice_l173_367;
  wire                when_ArraySlice_l285_6;
  wire                when_ArraySlice_l288_6;
  wire                outputStreamArrayData_6_fire_10;
  wire                when_ArraySlice_l292_6;
  wire                outputStreamArrayData_6_fire_11;
  wire                when_ArraySlice_l303_6;
  reg        [6:0]    _zz_when_ArraySlice_l304_6;
  wire       [5:0]    _zz_when_ArraySlice_l94_44;
  wire                when_ArraySlice_l94_44;
  wire                when_ArraySlice_l95_44;
  wire                when_ArraySlice_l99_44;
  wire                when_ArraySlice_l304_6;
  reg                 debug_0_46 /* verilator public */ ;
  reg                 debug_1_46 /* verilator public */ ;
  reg                 debug_2_46 /* verilator public */ ;
  reg                 debug_3_46 /* verilator public */ ;
  reg                 debug_4_46 /* verilator public */ ;
  reg                 debug_5_46 /* verilator public */ ;
  reg                 debug_6_46 /* verilator public */ ;
  reg                 debug_7_46 /* verilator public */ ;
  wire                when_ArraySlice_l165_368;
  wire                when_ArraySlice_l166_368;
  reg        [6:0]    _zz_when_ArraySlice_l173_368;
  wire       [5:0]    _zz_when_ArraySlice_l112_368;
  wire                when_ArraySlice_l112_368;
  wire                when_ArraySlice_l113_368;
  wire                when_ArraySlice_l118_368;
  wire                when_ArraySlice_l173_368;
  wire                when_ArraySlice_l165_369;
  wire                when_ArraySlice_l166_369;
  reg        [6:0]    _zz_when_ArraySlice_l173_369;
  wire       [5:0]    _zz_when_ArraySlice_l112_369;
  wire                when_ArraySlice_l112_369;
  wire                when_ArraySlice_l113_369;
  wire                when_ArraySlice_l118_369;
  wire                when_ArraySlice_l173_369;
  wire                when_ArraySlice_l165_370;
  wire                when_ArraySlice_l166_370;
  reg        [6:0]    _zz_when_ArraySlice_l173_370;
  wire       [5:0]    _zz_when_ArraySlice_l112_370;
  wire                when_ArraySlice_l112_370;
  wire                when_ArraySlice_l113_370;
  wire                when_ArraySlice_l118_370;
  wire                when_ArraySlice_l173_370;
  wire                when_ArraySlice_l165_371;
  wire                when_ArraySlice_l166_371;
  reg        [6:0]    _zz_when_ArraySlice_l173_371;
  wire       [5:0]    _zz_when_ArraySlice_l112_371;
  wire                when_ArraySlice_l112_371;
  wire                when_ArraySlice_l113_371;
  wire                when_ArraySlice_l118_371;
  wire                when_ArraySlice_l173_371;
  wire                when_ArraySlice_l165_372;
  wire                when_ArraySlice_l166_372;
  reg        [6:0]    _zz_when_ArraySlice_l173_372;
  wire       [5:0]    _zz_when_ArraySlice_l112_372;
  wire                when_ArraySlice_l112_372;
  wire                when_ArraySlice_l113_372;
  wire                when_ArraySlice_l118_372;
  wire                when_ArraySlice_l173_372;
  wire                when_ArraySlice_l165_373;
  wire                when_ArraySlice_l166_373;
  reg        [6:0]    _zz_when_ArraySlice_l173_373;
  wire       [5:0]    _zz_when_ArraySlice_l112_373;
  wire                when_ArraySlice_l112_373;
  wire                when_ArraySlice_l113_373;
  wire                when_ArraySlice_l118_373;
  wire                when_ArraySlice_l173_373;
  wire                when_ArraySlice_l165_374;
  wire                when_ArraySlice_l166_374;
  reg        [6:0]    _zz_when_ArraySlice_l173_374;
  wire       [5:0]    _zz_when_ArraySlice_l112_374;
  wire                when_ArraySlice_l112_374;
  wire                when_ArraySlice_l113_374;
  wire                when_ArraySlice_l118_374;
  wire                when_ArraySlice_l173_374;
  wire                when_ArraySlice_l165_375;
  wire                when_ArraySlice_l166_375;
  reg        [6:0]    _zz_when_ArraySlice_l173_375;
  wire       [5:0]    _zz_when_ArraySlice_l112_375;
  wire                when_ArraySlice_l112_375;
  wire                when_ArraySlice_l113_375;
  wire                when_ArraySlice_l118_375;
  wire                when_ArraySlice_l173_375;
  wire                when_ArraySlice_l311_6;
  wire                outputStreamArrayData_6_fire_12;
  wire                when_ArraySlice_l315_6;
  wire                when_ArraySlice_l301_6;
  wire                outputStreamArrayData_6_fire_13;
  wire                when_ArraySlice_l322_6;
  wire                when_ArraySlice_l240_7;
  wire                when_ArraySlice_l241_7;
  wire       [5:0]    _zz_outputStreamArrayData_7_valid_1;
  wire                _zz_io_pop_ready_15;
  wire       [63:0]   _zz_18;
  wire                when_ArraySlice_l246_7;
  wire                outputStreamArrayData_7_fire_7;
  wire                when_ArraySlice_l247_7;
  wire                when_ArraySlice_l248_7;
  wire                when_ArraySlice_l251_7;
  wire                outputStreamArrayData_7_fire_8;
  wire                when_ArraySlice_l256_7;
  wire                when_ArraySlice_l257_7;
  reg        [6:0]    _zz_when_ArraySlice_l259_7;
  wire       [5:0]    _zz_when_ArraySlice_l94_45;
  wire                when_ArraySlice_l94_45;
  wire                when_ArraySlice_l95_45;
  wire                when_ArraySlice_l99_45;
  wire                when_ArraySlice_l259_7;
  reg                 debug_0_47 /* verilator public */ ;
  reg                 debug_1_47 /* verilator public */ ;
  reg                 debug_2_47 /* verilator public */ ;
  reg                 debug_3_47 /* verilator public */ ;
  reg                 debug_4_47 /* verilator public */ ;
  reg                 debug_5_47 /* verilator public */ ;
  reg                 debug_6_47 /* verilator public */ ;
  reg                 debug_7_47 /* verilator public */ ;
  wire                when_ArraySlice_l165_376;
  wire                when_ArraySlice_l166_376;
  reg        [6:0]    _zz_when_ArraySlice_l173_376;
  wire       [5:0]    _zz_when_ArraySlice_l112_376;
  wire                when_ArraySlice_l112_376;
  wire                when_ArraySlice_l113_376;
  wire                when_ArraySlice_l118_376;
  wire                when_ArraySlice_l173_376;
  wire                when_ArraySlice_l165_377;
  wire                when_ArraySlice_l166_377;
  reg        [6:0]    _zz_when_ArraySlice_l173_377;
  wire       [5:0]    _zz_when_ArraySlice_l112_377;
  wire                when_ArraySlice_l112_377;
  wire                when_ArraySlice_l113_377;
  wire                when_ArraySlice_l118_377;
  wire                when_ArraySlice_l173_377;
  wire                when_ArraySlice_l165_378;
  wire                when_ArraySlice_l166_378;
  reg        [6:0]    _zz_when_ArraySlice_l173_378;
  wire       [5:0]    _zz_when_ArraySlice_l112_378;
  wire                when_ArraySlice_l112_378;
  wire                when_ArraySlice_l113_378;
  wire                when_ArraySlice_l118_378;
  wire                when_ArraySlice_l173_378;
  wire                when_ArraySlice_l165_379;
  wire                when_ArraySlice_l166_379;
  reg        [6:0]    _zz_when_ArraySlice_l173_379;
  wire       [5:0]    _zz_when_ArraySlice_l112_379;
  wire                when_ArraySlice_l112_379;
  wire                when_ArraySlice_l113_379;
  wire                when_ArraySlice_l118_379;
  wire                when_ArraySlice_l173_379;
  wire                when_ArraySlice_l165_380;
  wire                when_ArraySlice_l166_380;
  reg        [6:0]    _zz_when_ArraySlice_l173_380;
  wire       [5:0]    _zz_when_ArraySlice_l112_380;
  wire                when_ArraySlice_l112_380;
  wire                when_ArraySlice_l113_380;
  wire                when_ArraySlice_l118_380;
  wire                when_ArraySlice_l173_380;
  wire                when_ArraySlice_l165_381;
  wire                when_ArraySlice_l166_381;
  reg        [6:0]    _zz_when_ArraySlice_l173_381;
  wire       [5:0]    _zz_when_ArraySlice_l112_381;
  wire                when_ArraySlice_l112_381;
  wire                when_ArraySlice_l113_381;
  wire                when_ArraySlice_l118_381;
  wire                when_ArraySlice_l173_381;
  wire                when_ArraySlice_l165_382;
  wire                when_ArraySlice_l166_382;
  reg        [6:0]    _zz_when_ArraySlice_l173_382;
  wire       [5:0]    _zz_when_ArraySlice_l112_382;
  wire                when_ArraySlice_l112_382;
  wire                when_ArraySlice_l113_382;
  wire                when_ArraySlice_l118_382;
  wire                when_ArraySlice_l173_382;
  wire                when_ArraySlice_l165_383;
  wire                when_ArraySlice_l166_383;
  reg        [6:0]    _zz_when_ArraySlice_l173_383;
  wire       [5:0]    _zz_when_ArraySlice_l112_383;
  wire                when_ArraySlice_l112_383;
  wire                when_ArraySlice_l113_383;
  wire                when_ArraySlice_l118_383;
  wire                when_ArraySlice_l173_383;
  wire                when_ArraySlice_l265_7;
  wire                when_ArraySlice_l268_7;
  wire                when_ArraySlice_l272_7;
  wire                when_ArraySlice_l276_7;
  wire                outputStreamArrayData_7_fire_9;
  wire                when_ArraySlice_l277_7;
  reg        [6:0]    _zz_when_ArraySlice_l279_7;
  wire       [5:0]    _zz_when_ArraySlice_l94_46;
  wire                when_ArraySlice_l94_46;
  wire                when_ArraySlice_l95_46;
  wire                when_ArraySlice_l99_46;
  wire                when_ArraySlice_l279_7;
  reg                 debug_0_48 /* verilator public */ ;
  reg                 debug_1_48 /* verilator public */ ;
  reg                 debug_2_48 /* verilator public */ ;
  reg                 debug_3_48 /* verilator public */ ;
  reg                 debug_4_48 /* verilator public */ ;
  reg                 debug_5_48 /* verilator public */ ;
  reg                 debug_6_48 /* verilator public */ ;
  reg                 debug_7_48 /* verilator public */ ;
  wire                when_ArraySlice_l165_384;
  wire                when_ArraySlice_l166_384;
  reg        [6:0]    _zz_when_ArraySlice_l173_384;
  wire       [5:0]    _zz_when_ArraySlice_l112_384;
  wire                when_ArraySlice_l112_384;
  wire                when_ArraySlice_l113_384;
  wire                when_ArraySlice_l118_384;
  wire                when_ArraySlice_l173_384;
  wire                when_ArraySlice_l165_385;
  wire                when_ArraySlice_l166_385;
  reg        [6:0]    _zz_when_ArraySlice_l173_385;
  wire       [5:0]    _zz_when_ArraySlice_l112_385;
  wire                when_ArraySlice_l112_385;
  wire                when_ArraySlice_l113_385;
  wire                when_ArraySlice_l118_385;
  wire                when_ArraySlice_l173_385;
  wire                when_ArraySlice_l165_386;
  wire                when_ArraySlice_l166_386;
  reg        [6:0]    _zz_when_ArraySlice_l173_386;
  wire       [5:0]    _zz_when_ArraySlice_l112_386;
  wire                when_ArraySlice_l112_386;
  wire                when_ArraySlice_l113_386;
  wire                when_ArraySlice_l118_386;
  wire                when_ArraySlice_l173_386;
  wire                when_ArraySlice_l165_387;
  wire                when_ArraySlice_l166_387;
  reg        [6:0]    _zz_when_ArraySlice_l173_387;
  wire       [5:0]    _zz_when_ArraySlice_l112_387;
  wire                when_ArraySlice_l112_387;
  wire                when_ArraySlice_l113_387;
  wire                when_ArraySlice_l118_387;
  wire                when_ArraySlice_l173_387;
  wire                when_ArraySlice_l165_388;
  wire                when_ArraySlice_l166_388;
  reg        [6:0]    _zz_when_ArraySlice_l173_388;
  wire       [5:0]    _zz_when_ArraySlice_l112_388;
  wire                when_ArraySlice_l112_388;
  wire                when_ArraySlice_l113_388;
  wire                when_ArraySlice_l118_388;
  wire                when_ArraySlice_l173_388;
  wire                when_ArraySlice_l165_389;
  wire                when_ArraySlice_l166_389;
  reg        [6:0]    _zz_when_ArraySlice_l173_389;
  wire       [5:0]    _zz_when_ArraySlice_l112_389;
  wire                when_ArraySlice_l112_389;
  wire                when_ArraySlice_l113_389;
  wire                when_ArraySlice_l118_389;
  wire                when_ArraySlice_l173_389;
  wire                when_ArraySlice_l165_390;
  wire                when_ArraySlice_l166_390;
  reg        [6:0]    _zz_when_ArraySlice_l173_390;
  wire       [5:0]    _zz_when_ArraySlice_l112_390;
  wire                when_ArraySlice_l112_390;
  wire                when_ArraySlice_l113_390;
  wire                when_ArraySlice_l118_390;
  wire                when_ArraySlice_l173_390;
  wire                when_ArraySlice_l165_391;
  wire                when_ArraySlice_l166_391;
  reg        [6:0]    _zz_when_ArraySlice_l173_391;
  wire       [5:0]    _zz_when_ArraySlice_l112_391;
  wire                when_ArraySlice_l112_391;
  wire                when_ArraySlice_l113_391;
  wire                when_ArraySlice_l118_391;
  wire                when_ArraySlice_l173_391;
  wire                when_ArraySlice_l285_7;
  wire                when_ArraySlice_l288_7;
  wire                outputStreamArrayData_7_fire_10;
  wire                when_ArraySlice_l292_7;
  wire                outputStreamArrayData_7_fire_11;
  wire                when_ArraySlice_l303_7;
  reg        [6:0]    _zz_when_ArraySlice_l304_7;
  wire       [5:0]    _zz_when_ArraySlice_l94_47;
  wire                when_ArraySlice_l94_47;
  wire                when_ArraySlice_l95_47;
  wire                when_ArraySlice_l99_47;
  wire                when_ArraySlice_l304_7;
  reg                 debug_0_49 /* verilator public */ ;
  reg                 debug_1_49 /* verilator public */ ;
  reg                 debug_2_49 /* verilator public */ ;
  reg                 debug_3_49 /* verilator public */ ;
  reg                 debug_4_49 /* verilator public */ ;
  reg                 debug_5_49 /* verilator public */ ;
  reg                 debug_6_49 /* verilator public */ ;
  reg                 debug_7_49 /* verilator public */ ;
  wire                when_ArraySlice_l165_392;
  wire                when_ArraySlice_l166_392;
  reg        [6:0]    _zz_when_ArraySlice_l173_392;
  wire       [5:0]    _zz_when_ArraySlice_l112_392;
  wire                when_ArraySlice_l112_392;
  wire                when_ArraySlice_l113_392;
  wire                when_ArraySlice_l118_392;
  wire                when_ArraySlice_l173_392;
  wire                when_ArraySlice_l165_393;
  wire                when_ArraySlice_l166_393;
  reg        [6:0]    _zz_when_ArraySlice_l173_393;
  wire       [5:0]    _zz_when_ArraySlice_l112_393;
  wire                when_ArraySlice_l112_393;
  wire                when_ArraySlice_l113_393;
  wire                when_ArraySlice_l118_393;
  wire                when_ArraySlice_l173_393;
  wire                when_ArraySlice_l165_394;
  wire                when_ArraySlice_l166_394;
  reg        [6:0]    _zz_when_ArraySlice_l173_394;
  wire       [5:0]    _zz_when_ArraySlice_l112_394;
  wire                when_ArraySlice_l112_394;
  wire                when_ArraySlice_l113_394;
  wire                when_ArraySlice_l118_394;
  wire                when_ArraySlice_l173_394;
  wire                when_ArraySlice_l165_395;
  wire                when_ArraySlice_l166_395;
  reg        [6:0]    _zz_when_ArraySlice_l173_395;
  wire       [5:0]    _zz_when_ArraySlice_l112_395;
  wire                when_ArraySlice_l112_395;
  wire                when_ArraySlice_l113_395;
  wire                when_ArraySlice_l118_395;
  wire                when_ArraySlice_l173_395;
  wire                when_ArraySlice_l165_396;
  wire                when_ArraySlice_l166_396;
  reg        [6:0]    _zz_when_ArraySlice_l173_396;
  wire       [5:0]    _zz_when_ArraySlice_l112_396;
  wire                when_ArraySlice_l112_396;
  wire                when_ArraySlice_l113_396;
  wire                when_ArraySlice_l118_396;
  wire                when_ArraySlice_l173_396;
  wire                when_ArraySlice_l165_397;
  wire                when_ArraySlice_l166_397;
  reg        [6:0]    _zz_when_ArraySlice_l173_397;
  wire       [5:0]    _zz_when_ArraySlice_l112_397;
  wire                when_ArraySlice_l112_397;
  wire                when_ArraySlice_l113_397;
  wire                when_ArraySlice_l118_397;
  wire                when_ArraySlice_l173_397;
  wire                when_ArraySlice_l165_398;
  wire                when_ArraySlice_l166_398;
  reg        [6:0]    _zz_when_ArraySlice_l173_398;
  wire       [5:0]    _zz_when_ArraySlice_l112_398;
  wire                when_ArraySlice_l112_398;
  wire                when_ArraySlice_l113_398;
  wire                when_ArraySlice_l118_398;
  wire                when_ArraySlice_l173_398;
  wire                when_ArraySlice_l165_399;
  wire                when_ArraySlice_l166_399;
  reg        [6:0]    _zz_when_ArraySlice_l173_399;
  wire       [5:0]    _zz_when_ArraySlice_l112_399;
  wire                when_ArraySlice_l112_399;
  wire                when_ArraySlice_l113_399;
  wire                when_ArraySlice_l118_399;
  wire                when_ArraySlice_l173_399;
  wire                when_ArraySlice_l311_7;
  wire                outputStreamArrayData_7_fire_12;
  wire                when_ArraySlice_l315_7;
  wire                when_ArraySlice_l301_7;
  wire                outputStreamArrayData_7_fire_13;
  wire                when_ArraySlice_l322_7;
  reg                 _zz_when_ArraySlice_l333;
  reg                 _zz_when_ArraySlice_l333_1;
  reg                 _zz_when_ArraySlice_l333_2;
  reg                 _zz_when_ArraySlice_l333_3;
  reg                 _zz_when_ArraySlice_l333_4;
  reg                 _zz_when_ArraySlice_l333_5;
  reg                 _zz_when_ArraySlice_l333_6;
  reg                 _zz_when_ArraySlice_l333_7;
  wire                when_ArraySlice_l189;
  wire                when_ArraySlice_l190;
  wire                when_ArraySlice_l189_1;
  wire                when_ArraySlice_l190_1;
  wire                when_ArraySlice_l189_2;
  wire                when_ArraySlice_l190_2;
  wire                when_ArraySlice_l189_3;
  wire                when_ArraySlice_l190_3;
  wire                when_ArraySlice_l189_4;
  wire                when_ArraySlice_l190_4;
  wire                when_ArraySlice_l189_5;
  wire                when_ArraySlice_l190_5;
  wire                when_ArraySlice_l189_6;
  wire                when_ArraySlice_l190_6;
  wire                when_ArraySlice_l189_7;
  wire                when_ArraySlice_l190_7;
  wire                when_ArraySlice_l333;
  wire                when_ArraySlice_l334;
  wire                _zz_io_push_valid_1;
  wire       [31:0]   _zz_io_push_payload_1;
  wire       [63:0]   _zz_19;
  wire       [63:0]   _zz_20;
  wire                inputStreamArrayData_fire_1;
  wire                when_ArraySlice_l338;
  wire                when_ArraySlice_l339;
  reg                 debug_0_50 /* verilator public */ ;
  reg                 debug_1_50 /* verilator public */ ;
  reg                 debug_2_50 /* verilator public */ ;
  reg                 debug_3_50 /* verilator public */ ;
  reg                 debug_4_50 /* verilator public */ ;
  reg                 debug_5_50 /* verilator public */ ;
  reg                 debug_6_50 /* verilator public */ ;
  reg                 debug_7_50 /* verilator public */ ;
  wire                when_ArraySlice_l165_400;
  wire                when_ArraySlice_l166_400;
  reg        [6:0]    _zz_when_ArraySlice_l173_400;
  wire       [5:0]    _zz_when_ArraySlice_l112_400;
  wire                when_ArraySlice_l112_400;
  wire                when_ArraySlice_l113_400;
  wire                when_ArraySlice_l118_400;
  wire                when_ArraySlice_l173_400;
  wire                when_ArraySlice_l165_401;
  wire                when_ArraySlice_l166_401;
  reg        [6:0]    _zz_when_ArraySlice_l173_401;
  wire       [5:0]    _zz_when_ArraySlice_l112_401;
  wire                when_ArraySlice_l112_401;
  wire                when_ArraySlice_l113_401;
  wire                when_ArraySlice_l118_401;
  wire                when_ArraySlice_l173_401;
  wire                when_ArraySlice_l165_402;
  wire                when_ArraySlice_l166_402;
  reg        [6:0]    _zz_when_ArraySlice_l173_402;
  wire       [5:0]    _zz_when_ArraySlice_l112_402;
  wire                when_ArraySlice_l112_402;
  wire                when_ArraySlice_l113_402;
  wire                when_ArraySlice_l118_402;
  wire                when_ArraySlice_l173_402;
  wire                when_ArraySlice_l165_403;
  wire                when_ArraySlice_l166_403;
  reg        [6:0]    _zz_when_ArraySlice_l173_403;
  wire       [5:0]    _zz_when_ArraySlice_l112_403;
  wire                when_ArraySlice_l112_403;
  wire                when_ArraySlice_l113_403;
  wire                when_ArraySlice_l118_403;
  wire                when_ArraySlice_l173_403;
  wire                when_ArraySlice_l165_404;
  wire                when_ArraySlice_l166_404;
  reg        [6:0]    _zz_when_ArraySlice_l173_404;
  wire       [5:0]    _zz_when_ArraySlice_l112_404;
  wire                when_ArraySlice_l112_404;
  wire                when_ArraySlice_l113_404;
  wire                when_ArraySlice_l118_404;
  wire                when_ArraySlice_l173_404;
  wire                when_ArraySlice_l165_405;
  wire                when_ArraySlice_l166_405;
  reg        [6:0]    _zz_when_ArraySlice_l173_405;
  wire       [5:0]    _zz_when_ArraySlice_l112_405;
  wire                when_ArraySlice_l112_405;
  wire                when_ArraySlice_l113_405;
  wire                when_ArraySlice_l118_405;
  wire                when_ArraySlice_l173_405;
  wire                when_ArraySlice_l165_406;
  wire                when_ArraySlice_l166_406;
  reg        [6:0]    _zz_when_ArraySlice_l173_406;
  wire       [5:0]    _zz_when_ArraySlice_l112_406;
  wire                when_ArraySlice_l112_406;
  wire                when_ArraySlice_l113_406;
  wire                when_ArraySlice_l118_406;
  wire                when_ArraySlice_l173_406;
  wire                when_ArraySlice_l165_407;
  wire                when_ArraySlice_l166_407;
  reg        [6:0]    _zz_when_ArraySlice_l173_407;
  wire       [5:0]    _zz_when_ArraySlice_l112_407;
  wire                when_ArraySlice_l112_407;
  wire                when_ArraySlice_l113_407;
  wire                when_ArraySlice_l118_407;
  wire                when_ArraySlice_l173_407;
  wire                when_ArraySlice_l350;
  reg                 debug_0_51 /* verilator public */ ;
  reg                 debug_1_51 /* verilator public */ ;
  reg                 debug_2_51 /* verilator public */ ;
  reg                 debug_3_51 /* verilator public */ ;
  reg                 debug_4_51 /* verilator public */ ;
  reg                 debug_5_51 /* verilator public */ ;
  reg                 debug_6_51 /* verilator public */ ;
  reg                 debug_7_51 /* verilator public */ ;
  wire                when_ArraySlice_l165_408;
  wire                when_ArraySlice_l166_408;
  reg        [6:0]    _zz_when_ArraySlice_l173_408;
  wire       [5:0]    _zz_when_ArraySlice_l112_408;
  wire                when_ArraySlice_l112_408;
  wire                when_ArraySlice_l113_408;
  wire                when_ArraySlice_l118_408;
  wire                when_ArraySlice_l173_408;
  wire                when_ArraySlice_l165_409;
  wire                when_ArraySlice_l166_409;
  reg        [6:0]    _zz_when_ArraySlice_l173_409;
  wire       [5:0]    _zz_when_ArraySlice_l112_409;
  wire                when_ArraySlice_l112_409;
  wire                when_ArraySlice_l113_409;
  wire                when_ArraySlice_l118_409;
  wire                when_ArraySlice_l173_409;
  wire                when_ArraySlice_l165_410;
  wire                when_ArraySlice_l166_410;
  reg        [6:0]    _zz_when_ArraySlice_l173_410;
  wire       [5:0]    _zz_when_ArraySlice_l112_410;
  wire                when_ArraySlice_l112_410;
  wire                when_ArraySlice_l113_410;
  wire                when_ArraySlice_l118_410;
  wire                when_ArraySlice_l173_410;
  wire                when_ArraySlice_l165_411;
  wire                when_ArraySlice_l166_411;
  reg        [6:0]    _zz_when_ArraySlice_l173_411;
  wire       [5:0]    _zz_when_ArraySlice_l112_411;
  wire                when_ArraySlice_l112_411;
  wire                when_ArraySlice_l113_411;
  wire                when_ArraySlice_l118_411;
  wire                when_ArraySlice_l173_411;
  wire                when_ArraySlice_l165_412;
  wire                when_ArraySlice_l166_412;
  reg        [6:0]    _zz_when_ArraySlice_l173_412;
  wire       [5:0]    _zz_when_ArraySlice_l112_412;
  wire                when_ArraySlice_l112_412;
  wire                when_ArraySlice_l113_412;
  wire                when_ArraySlice_l118_412;
  wire                when_ArraySlice_l173_412;
  wire                when_ArraySlice_l165_413;
  wire                when_ArraySlice_l166_413;
  reg        [6:0]    _zz_when_ArraySlice_l173_413;
  wire       [5:0]    _zz_when_ArraySlice_l112_413;
  wire                when_ArraySlice_l112_413;
  wire                when_ArraySlice_l113_413;
  wire                when_ArraySlice_l118_413;
  wire                when_ArraySlice_l173_413;
  wire                when_ArraySlice_l165_414;
  wire                when_ArraySlice_l166_414;
  reg        [6:0]    _zz_when_ArraySlice_l173_414;
  wire       [5:0]    _zz_when_ArraySlice_l112_414;
  wire                when_ArraySlice_l112_414;
  wire                when_ArraySlice_l113_414;
  wire                when_ArraySlice_l118_414;
  wire                when_ArraySlice_l173_414;
  wire                when_ArraySlice_l165_415;
  wire                when_ArraySlice_l166_415;
  reg        [6:0]    _zz_when_ArraySlice_l173_415;
  wire       [5:0]    _zz_when_ArraySlice_l112_415;
  wire                when_ArraySlice_l112_415;
  wire                when_ArraySlice_l113_415;
  wire                when_ArraySlice_l118_415;
  wire                when_ArraySlice_l173_415;
  reg                 _zz_when_ArraySlice_l354;
  reg                 _zz_when_ArraySlice_l354_1;
  reg                 _zz_when_ArraySlice_l354_2;
  reg                 _zz_when_ArraySlice_l354_3;
  reg                 _zz_when_ArraySlice_l354_4;
  reg                 _zz_when_ArraySlice_l354_5;
  reg                 _zz_when_ArraySlice_l354_6;
  reg                 _zz_when_ArraySlice_l354_7;
  wire                when_ArraySlice_l189_8;
  wire                when_ArraySlice_l190_8;
  wire                when_ArraySlice_l189_9;
  wire                when_ArraySlice_l190_9;
  wire                when_ArraySlice_l189_10;
  wire                when_ArraySlice_l190_10;
  wire                when_ArraySlice_l189_11;
  wire                when_ArraySlice_l190_11;
  wire                when_ArraySlice_l189_12;
  wire                when_ArraySlice_l190_12;
  wire                when_ArraySlice_l189_13;
  wire                when_ArraySlice_l190_13;
  wire                when_ArraySlice_l189_14;
  wire                when_ArraySlice_l190_14;
  wire                when_ArraySlice_l189_15;
  wire                when_ArraySlice_l190_15;
  wire                when_ArraySlice_l354;
  reg                 _zz_when_ArraySlice_l358;
  reg                 _zz_when_ArraySlice_l358_1;
  reg                 _zz_when_ArraySlice_l358_2;
  reg                 _zz_when_ArraySlice_l358_3;
  reg                 _zz_when_ArraySlice_l358_4;
  reg                 _zz_when_ArraySlice_l358_5;
  reg                 _zz_when_ArraySlice_l358_6;
  reg                 _zz_when_ArraySlice_l358_7;
  wire                when_ArraySlice_l189_16;
  wire                when_ArraySlice_l190_16;
  wire                when_ArraySlice_l189_17;
  wire                when_ArraySlice_l190_17;
  wire                when_ArraySlice_l189_18;
  wire                when_ArraySlice_l190_18;
  wire                when_ArraySlice_l189_19;
  wire                when_ArraySlice_l190_19;
  wire                when_ArraySlice_l189_20;
  wire                when_ArraySlice_l190_20;
  wire                when_ArraySlice_l189_21;
  wire                when_ArraySlice_l190_21;
  wire                when_ArraySlice_l189_22;
  wire                when_ArraySlice_l190_22;
  wire                when_ArraySlice_l189_23;
  wire                when_ArraySlice_l190_23;
  wire                when_ArraySlice_l358;
  wire                when_ArraySlice_l361;
  wire                when_ArraySlice_l361_1;
  wire                when_ArraySlice_l361_2;
  wire                when_ArraySlice_l361_3;
  wire                when_ArraySlice_l361_4;
  wire                when_ArraySlice_l361_5;
  wire                when_ArraySlice_l361_6;
  wire                when_ArraySlice_l361_7;
  `ifndef SYNTHESIS
  reg [103:0] arraySliceStateMachine_stateReg_string;
  reg [103:0] arraySliceStateMachine_stateNext_string;
  `endif


  assign _zz_handshakeTimes_0_valueNext_1 = handshakeTimes_0_willIncrement;
  assign _zz_handshakeTimes_0_valueNext = {12'd0, _zz_handshakeTimes_0_valueNext_1};
  assign _zz_handshakeTimes_1_valueNext_1 = handshakeTimes_1_willIncrement;
  assign _zz_handshakeTimes_1_valueNext = {12'd0, _zz_handshakeTimes_1_valueNext_1};
  assign _zz_handshakeTimes_2_valueNext_1 = handshakeTimes_2_willIncrement;
  assign _zz_handshakeTimes_2_valueNext = {12'd0, _zz_handshakeTimes_2_valueNext_1};
  assign _zz_handshakeTimes_3_valueNext_1 = handshakeTimes_3_willIncrement;
  assign _zz_handshakeTimes_3_valueNext = {12'd0, _zz_handshakeTimes_3_valueNext_1};
  assign _zz_handshakeTimes_4_valueNext_1 = handshakeTimes_4_willIncrement;
  assign _zz_handshakeTimes_4_valueNext = {12'd0, _zz_handshakeTimes_4_valueNext_1};
  assign _zz_handshakeTimes_5_valueNext_1 = handshakeTimes_5_willIncrement;
  assign _zz_handshakeTimes_5_valueNext = {12'd0, _zz_handshakeTimes_5_valueNext_1};
  assign _zz_handshakeTimes_6_valueNext_1 = handshakeTimes_6_willIncrement;
  assign _zz_handshakeTimes_6_valueNext = {12'd0, _zz_handshakeTimes_6_valueNext_1};
  assign _zz_handshakeTimes_7_valueNext_1 = handshakeTimes_7_willIncrement;
  assign _zz_handshakeTimes_7_valueNext = {12'd0, _zz_handshakeTimes_7_valueNext_1};
  assign _zz_outSliceNumb_0_valueNext_1 = outSliceNumb_0_willIncrement;
  assign _zz_outSliceNumb_0_valueNext = {6'd0, _zz_outSliceNumb_0_valueNext_1};
  assign _zz_outSliceNumb_1_valueNext_1 = outSliceNumb_1_willIncrement;
  assign _zz_outSliceNumb_1_valueNext = {6'd0, _zz_outSliceNumb_1_valueNext_1};
  assign _zz_outSliceNumb_2_valueNext_1 = outSliceNumb_2_willIncrement;
  assign _zz_outSliceNumb_2_valueNext = {6'd0, _zz_outSliceNumb_2_valueNext_1};
  assign _zz_outSliceNumb_3_valueNext_1 = outSliceNumb_3_willIncrement;
  assign _zz_outSliceNumb_3_valueNext = {6'd0, _zz_outSliceNumb_3_valueNext_1};
  assign _zz_outSliceNumb_4_valueNext_1 = outSliceNumb_4_willIncrement;
  assign _zz_outSliceNumb_4_valueNext = {6'd0, _zz_outSliceNumb_4_valueNext_1};
  assign _zz_outSliceNumb_5_valueNext_1 = outSliceNumb_5_willIncrement;
  assign _zz_outSliceNumb_5_valueNext = {6'd0, _zz_outSliceNumb_5_valueNext_1};
  assign _zz_outSliceNumb_6_valueNext_1 = outSliceNumb_6_willIncrement;
  assign _zz_outSliceNumb_6_valueNext = {6'd0, _zz_outSliceNumb_6_valueNext_1};
  assign _zz_outSliceNumb_7_valueNext_1 = outSliceNumb_7_willIncrement;
  assign _zz_outSliceNumb_7_valueNext = {6'd0, _zz_outSliceNumb_7_valueNext_1};
  assign _zz_when_ArraySlice_l211_1 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l215_2 = (hReg - _zz_when_ArraySlice_l215_3);
  assign _zz_when_ArraySlice_l215_1 = {1'd0, _zz_when_ArraySlice_l215_2};
  assign _zz_when_ArraySlice_l215_4 = 1'b1;
  assign _zz_when_ArraySlice_l215_3 = {5'd0, _zz_when_ArraySlice_l215_4};
  assign _zz_when_ArraySlice_l216 = (wReg - _zz_when_ArraySlice_l216_1);
  assign _zz_when_ArraySlice_l216_2 = 1'b1;
  assign _zz_when_ArraySlice_l216_1 = {5'd0, _zz_when_ArraySlice_l216_2};
  assign _zz_selectWriteFifo_1 = 1'b1;
  assign _zz_selectWriteFifo = {5'd0, _zz_selectWriteFifo_1};
  assign _zz_when_ArraySlice_l165 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_1);
  assign _zz_when_ArraySlice_l165_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_1 = {3'd0, _zz_when_ArraySlice_l165_2};
  assign _zz_when_ArraySlice_l166 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_3);
  assign _zz_when_ArraySlice_l166_1 = {1'd0, _zz_when_ArraySlice_l166_2};
  assign _zz_when_ArraySlice_l166_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_4);
  assign _zz_when_ArraySlice_l166_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_4 = {3'd0, _zz_when_ArraySlice_l166_5};
  assign _zz__zz_when_ArraySlice_l112 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113 = (_zz_when_ArraySlice_l113_1 - _zz_when_ArraySlice_l113_4);
  assign _zz_when_ArraySlice_l113_1 = (_zz_when_ArraySlice_l113_2 + _zz_when_ArraySlice_l113_3);
  assign _zz_when_ArraySlice_l113_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_4 = {1'd0, _zz_when_ArraySlice_l112};
  assign _zz__zz_when_ArraySlice_l173 = (_zz__zz_when_ArraySlice_l173_1 + _zz__zz_when_ArraySlice_l173_2);
  assign _zz__zz_when_ArraySlice_l173_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_3 = {1'd0, _zz_when_ArraySlice_l112};
  assign _zz_when_ArraySlice_l118_1 = 7'h40;
  assign _zz_when_ArraySlice_l118 = _zz_when_ArraySlice_l118_1[5:0];
  assign _zz_when_ArraySlice_l173_416 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_417 = (_zz_when_ArraySlice_l173_418 + _zz_when_ArraySlice_l173_423);
  assign _zz_when_ArraySlice_l173_418 = (_zz_when_ArraySlice_l173 - _zz_when_ArraySlice_l173_419);
  assign _zz_when_ArraySlice_l173_420 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_421);
  assign _zz_when_ArraySlice_l173_419 = {1'd0, _zz_when_ArraySlice_l173_420};
  assign _zz_when_ArraySlice_l173_422 = 3'b000;
  assign _zz_when_ArraySlice_l173_421 = {3'd0, _zz_when_ArraySlice_l173_422};
  assign _zz_when_ArraySlice_l173_423 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_1_1 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_1_2);
  assign _zz_when_ArraySlice_l165_1_3 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_1_2 = {2'd0, _zz_when_ArraySlice_l165_1_3};
  assign _zz_when_ArraySlice_l166_1_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_1_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_1_3);
  assign _zz_when_ArraySlice_l166_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_1_4);
  assign _zz_when_ArraySlice_l166_1_5 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_1_4 = {2'd0, _zz_when_ArraySlice_l166_1_5};
  assign _zz__zz_when_ArraySlice_l112_1 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_1_1 = (_zz_when_ArraySlice_l113_1_2 - _zz_when_ArraySlice_l113_1_5);
  assign _zz_when_ArraySlice_l113_1_2 = (_zz_when_ArraySlice_l113_1_3 + _zz_when_ArraySlice_l113_1_4);
  assign _zz_when_ArraySlice_l113_1_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_1_4 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_1_5 = {1'd0, _zz_when_ArraySlice_l112_1};
  assign _zz__zz_when_ArraySlice_l173_1_1 = (_zz__zz_when_ArraySlice_l173_1_2 + _zz__zz_when_ArraySlice_l173_1_3);
  assign _zz__zz_when_ArraySlice_l173_1_2 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_1_3 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_1_4 = {1'd0, _zz_when_ArraySlice_l112_1};
  assign _zz_when_ArraySlice_l118_1_2 = 7'h40;
  assign _zz_when_ArraySlice_l118_1_1 = _zz_when_ArraySlice_l118_1_2[5:0];
  assign _zz_when_ArraySlice_l173_1_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_1_1 = {1'd0, _zz_when_ArraySlice_l173_1_2};
  assign _zz_when_ArraySlice_l173_1_3 = (_zz_when_ArraySlice_l173_1_4 + _zz_when_ArraySlice_l173_1_9);
  assign _zz_when_ArraySlice_l173_1_4 = (_zz_when_ArraySlice_l173_1 - _zz_when_ArraySlice_l173_1_5);
  assign _zz_when_ArraySlice_l173_1_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_1_7);
  assign _zz_when_ArraySlice_l173_1_5 = {1'd0, _zz_when_ArraySlice_l173_1_6};
  assign _zz_when_ArraySlice_l173_1_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_1_7 = {2'd0, _zz_when_ArraySlice_l173_1_8};
  assign _zz_when_ArraySlice_l173_1_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_2_1 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_2_2);
  assign _zz_when_ArraySlice_l165_2_3 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_2_2 = {1'd0, _zz_when_ArraySlice_l165_2_3};
  assign _zz_when_ArraySlice_l166_2_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_2_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_2_3);
  assign _zz_when_ArraySlice_l166_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_2_4);
  assign _zz_when_ArraySlice_l166_2_5 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_2_4 = {1'd0, _zz_when_ArraySlice_l166_2_5};
  assign _zz__zz_when_ArraySlice_l112_2 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_2_1 = (_zz_when_ArraySlice_l113_2_2 - _zz_when_ArraySlice_l113_2_5);
  assign _zz_when_ArraySlice_l113_2_2 = (_zz_when_ArraySlice_l113_2_3 + _zz_when_ArraySlice_l113_2_4);
  assign _zz_when_ArraySlice_l113_2_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_2_4 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_2_5 = {1'd0, _zz_when_ArraySlice_l112_2};
  assign _zz__zz_when_ArraySlice_l173_2_1 = (_zz__zz_when_ArraySlice_l173_2_2 + _zz__zz_when_ArraySlice_l173_2_3);
  assign _zz__zz_when_ArraySlice_l173_2_2 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_2_3 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_2_4 = {1'd0, _zz_when_ArraySlice_l112_2};
  assign _zz_when_ArraySlice_l118_2_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_2 = _zz_when_ArraySlice_l118_2_1[5:0];
  assign _zz_when_ArraySlice_l173_2_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_2_1 = {1'd0, _zz_when_ArraySlice_l173_2_2};
  assign _zz_when_ArraySlice_l173_2_3 = (_zz_when_ArraySlice_l173_2_4 + _zz_when_ArraySlice_l173_2_9);
  assign _zz_when_ArraySlice_l173_2_4 = (_zz_when_ArraySlice_l173_2 - _zz_when_ArraySlice_l173_2_5);
  assign _zz_when_ArraySlice_l173_2_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_2_7);
  assign _zz_when_ArraySlice_l173_2_5 = {1'd0, _zz_when_ArraySlice_l173_2_6};
  assign _zz_when_ArraySlice_l173_2_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_2_7 = {1'd0, _zz_when_ArraySlice_l173_2_8};
  assign _zz_when_ArraySlice_l173_2_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_3_1);
  assign _zz_when_ArraySlice_l165_3_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_3_1 = {1'd0, _zz_when_ArraySlice_l165_3_2};
  assign _zz_when_ArraySlice_l166_3_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_3_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_3_3);
  assign _zz_when_ArraySlice_l166_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_3_4);
  assign _zz_when_ArraySlice_l166_3_5 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_3_4 = {1'd0, _zz_when_ArraySlice_l166_3_5};
  assign _zz__zz_when_ArraySlice_l112_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_3_1 = (_zz_when_ArraySlice_l113_3_2 - _zz_when_ArraySlice_l113_3_5);
  assign _zz_when_ArraySlice_l113_3_2 = (_zz_when_ArraySlice_l113_3_3 + _zz_when_ArraySlice_l113_3_4);
  assign _zz_when_ArraySlice_l113_3_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_3_4 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_3_5 = {1'd0, _zz_when_ArraySlice_l112_3};
  assign _zz__zz_when_ArraySlice_l173_3_1 = (_zz__zz_when_ArraySlice_l173_3_2 + _zz__zz_when_ArraySlice_l173_3_3);
  assign _zz__zz_when_ArraySlice_l173_3_2 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_3_3 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_3_4 = {1'd0, _zz_when_ArraySlice_l112_3};
  assign _zz_when_ArraySlice_l118_3_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_3 = _zz_when_ArraySlice_l118_3_1[5:0];
  assign _zz_when_ArraySlice_l173_3_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_3_1 = {1'd0, _zz_when_ArraySlice_l173_3_2};
  assign _zz_when_ArraySlice_l173_3_3 = (_zz_when_ArraySlice_l173_3_4 + _zz_when_ArraySlice_l173_3_9);
  assign _zz_when_ArraySlice_l173_3_4 = (_zz_when_ArraySlice_l173_3 - _zz_when_ArraySlice_l173_3_5);
  assign _zz_when_ArraySlice_l173_3_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_3_7);
  assign _zz_when_ArraySlice_l173_3_5 = {1'd0, _zz_when_ArraySlice_l173_3_6};
  assign _zz_when_ArraySlice_l173_3_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_3_7 = {1'd0, _zz_when_ArraySlice_l173_3_8};
  assign _zz_when_ArraySlice_l173_3_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_4_1);
  assign _zz_when_ArraySlice_l165_4_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_4_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_4_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_4_3);
  assign _zz_when_ArraySlice_l166_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_4_4);
  assign _zz_when_ArraySlice_l166_4_4 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_4 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_4_1 = (_zz_when_ArraySlice_l113_4_2 - _zz_when_ArraySlice_l113_4_5);
  assign _zz_when_ArraySlice_l113_4_2 = (_zz_when_ArraySlice_l113_4_3 + _zz_when_ArraySlice_l113_4_4);
  assign _zz_when_ArraySlice_l113_4_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_4_4 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_4_5 = {1'd0, _zz_when_ArraySlice_l112_4};
  assign _zz__zz_when_ArraySlice_l173_4 = (_zz__zz_when_ArraySlice_l173_4_1 + _zz__zz_when_ArraySlice_l173_4_2);
  assign _zz__zz_when_ArraySlice_l173_4_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_4_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_4_3 = {1'd0, _zz_when_ArraySlice_l112_4};
  assign _zz_when_ArraySlice_l118_4_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_4 = _zz_when_ArraySlice_l118_4_1[5:0];
  assign _zz_when_ArraySlice_l173_4_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_4_1 = {1'd0, _zz_when_ArraySlice_l173_4_2};
  assign _zz_when_ArraySlice_l173_4_3 = (_zz_when_ArraySlice_l173_4_4 + _zz_when_ArraySlice_l173_4_8);
  assign _zz_when_ArraySlice_l173_4_4 = (_zz_when_ArraySlice_l173_4 - _zz_when_ArraySlice_l173_4_5);
  assign _zz_when_ArraySlice_l173_4_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_4_7);
  assign _zz_when_ArraySlice_l173_4_5 = {1'd0, _zz_when_ArraySlice_l173_4_6};
  assign _zz_when_ArraySlice_l173_4_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_4_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_5 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_5_1);
  assign _zz_when_ArraySlice_l165_5_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_5_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_5_1 = {1'd0, _zz_when_ArraySlice_l166_5_2};
  assign _zz_when_ArraySlice_l166_5_3 = (selectWriteFifo - _zz_when_ArraySlice_l166_5_4);
  assign _zz_when_ArraySlice_l166_5_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_5_5);
  assign _zz_when_ArraySlice_l166_5_5 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_5 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_5 = (_zz_when_ArraySlice_l113_5_1 - _zz_when_ArraySlice_l113_5_4);
  assign _zz_when_ArraySlice_l113_5_1 = (_zz_when_ArraySlice_l113_5_2 + _zz_when_ArraySlice_l113_5_3);
  assign _zz_when_ArraySlice_l113_5_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_5_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_5_4 = {1'd0, _zz_when_ArraySlice_l112_5};
  assign _zz__zz_when_ArraySlice_l173_5 = (_zz__zz_when_ArraySlice_l173_5_1 + _zz__zz_when_ArraySlice_l173_5_2);
  assign _zz__zz_when_ArraySlice_l173_5_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_5_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_5_3 = {1'd0, _zz_when_ArraySlice_l112_5};
  assign _zz_when_ArraySlice_l118_5_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_5 = _zz_when_ArraySlice_l118_5_1[5:0];
  assign _zz_when_ArraySlice_l173_5_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_5_1 = {2'd0, _zz_when_ArraySlice_l173_5_2};
  assign _zz_when_ArraySlice_l173_5_3 = (_zz_when_ArraySlice_l173_5_4 + _zz_when_ArraySlice_l173_5_8);
  assign _zz_when_ArraySlice_l173_5_4 = (_zz_when_ArraySlice_l173_5 - _zz_when_ArraySlice_l173_5_5);
  assign _zz_when_ArraySlice_l173_5_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_5_7);
  assign _zz_when_ArraySlice_l173_5_5 = {1'd0, _zz_when_ArraySlice_l173_5_6};
  assign _zz_when_ArraySlice_l173_5_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_5_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_6_1);
  assign _zz_when_ArraySlice_l165_6_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_6_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_6 = {1'd0, _zz_when_ArraySlice_l166_6_1};
  assign _zz_when_ArraySlice_l166_6_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_6_3);
  assign _zz_when_ArraySlice_l166_6_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_6_4);
  assign _zz_when_ArraySlice_l166_6_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_6 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_6 = (_zz_when_ArraySlice_l113_6_1 - _zz_when_ArraySlice_l113_6_4);
  assign _zz_when_ArraySlice_l113_6_1 = (_zz_when_ArraySlice_l113_6_2 + _zz_when_ArraySlice_l113_6_3);
  assign _zz_when_ArraySlice_l113_6_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_6_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_6_4 = {1'd0, _zz_when_ArraySlice_l112_6};
  assign _zz__zz_when_ArraySlice_l173_6 = (_zz__zz_when_ArraySlice_l173_6_1 + _zz__zz_when_ArraySlice_l173_6_2);
  assign _zz__zz_when_ArraySlice_l173_6_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_6_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_6_3 = {1'd0, _zz_when_ArraySlice_l112_6};
  assign _zz_when_ArraySlice_l118_6_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_6 = _zz_when_ArraySlice_l118_6_1[5:0];
  assign _zz_when_ArraySlice_l173_6_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_6_1 = {2'd0, _zz_when_ArraySlice_l173_6_2};
  assign _zz_when_ArraySlice_l173_6_3 = (_zz_when_ArraySlice_l173_6_4 + _zz_when_ArraySlice_l173_6_8);
  assign _zz_when_ArraySlice_l173_6_4 = (_zz_when_ArraySlice_l173_6 - _zz_when_ArraySlice_l173_6_5);
  assign _zz_when_ArraySlice_l173_6_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_6_7);
  assign _zz_when_ArraySlice_l173_6_5 = {1'd0, _zz_when_ArraySlice_l173_6_6};
  assign _zz_when_ArraySlice_l173_6_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_6_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_7 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_7_1);
  assign _zz_when_ArraySlice_l165_7_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_7_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_7 = {2'd0, _zz_when_ArraySlice_l166_7_1};
  assign _zz_when_ArraySlice_l166_7_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_7_3);
  assign _zz_when_ArraySlice_l166_7_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_7_4);
  assign _zz_when_ArraySlice_l166_7_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_7 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_7 = (_zz_when_ArraySlice_l113_7_1 - _zz_when_ArraySlice_l113_7_4);
  assign _zz_when_ArraySlice_l113_7_1 = (_zz_when_ArraySlice_l113_7_2 + _zz_when_ArraySlice_l113_7_3);
  assign _zz_when_ArraySlice_l113_7_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_7_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_7_4 = {1'd0, _zz_when_ArraySlice_l112_7};
  assign _zz__zz_when_ArraySlice_l173_7 = (_zz__zz_when_ArraySlice_l173_7_1 + _zz__zz_when_ArraySlice_l173_7_2);
  assign _zz__zz_when_ArraySlice_l173_7_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_7_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_7_3 = {1'd0, _zz_when_ArraySlice_l112_7};
  assign _zz_when_ArraySlice_l118_7_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_7 = _zz_when_ArraySlice_l118_7_1[5:0];
  assign _zz_when_ArraySlice_l173_7_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_7_1 = {3'd0, _zz_when_ArraySlice_l173_7_2};
  assign _zz_when_ArraySlice_l173_7_3 = (_zz_when_ArraySlice_l173_7_4 + _zz_when_ArraySlice_l173_7_8);
  assign _zz_when_ArraySlice_l173_7_4 = (_zz_when_ArraySlice_l173_7 - _zz_when_ArraySlice_l173_7_5);
  assign _zz_when_ArraySlice_l173_7_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_7_7);
  assign _zz_when_ArraySlice_l173_7_5 = {1'd0, _zz_when_ArraySlice_l173_7_6};
  assign _zz_when_ArraySlice_l173_7_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_7_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l373 = (selectReadFifo_0 + _zz_when_ArraySlice_l373_1);
  assign _zz_when_ArraySlice_l373_2 = 3'b000;
  assign _zz_when_ArraySlice_l373_1 = {3'd0, _zz_when_ArraySlice_l373_2};
  assign _zz_when_ArraySlice_l374_1 = (selectReadFifo_0 + _zz_when_ArraySlice_l374_2);
  assign _zz_when_ArraySlice_l374_3 = 3'b000;
  assign _zz_when_ArraySlice_l374_2 = {3'd0, _zz_when_ArraySlice_l374_3};
  assign _zz__zz_outputStreamArrayData_0_valid_1 = 3'b000;
  assign _zz__zz_outputStreamArrayData_0_valid = {3'd0, _zz__zz_outputStreamArrayData_0_valid_1};
  assign _zz_when_ArraySlice_l380_1 = 1'b1;
  assign _zz_when_ArraySlice_l380 = {6'd0, _zz_when_ArraySlice_l380_1};
  assign _zz_when_ArraySlice_l380_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l380_4);
  assign _zz_when_ArraySlice_l380_5 = 3'b000;
  assign _zz_when_ArraySlice_l380_4 = {3'd0, _zz_when_ArraySlice_l380_5};
  assign _zz_when_ArraySlice_l381_1 = (_zz_when_ArraySlice_l381_2 - _zz_when_ArraySlice_l381_3);
  assign _zz_when_ArraySlice_l381 = {7'd0, _zz_when_ArraySlice_l381_1};
  assign _zz_when_ArraySlice_l381_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l381_4 = 1'b1;
  assign _zz_when_ArraySlice_l381_3 = {5'd0, _zz_when_ArraySlice_l381_4};
  assign _zz_selectReadFifo_0 = (selectReadFifo_0 - _zz_selectReadFifo_0_1);
  assign _zz_selectReadFifo_0_1 = {3'd0, bReg};
  assign _zz_selectReadFifo_0_3 = 1'b1;
  assign _zz_selectReadFifo_0_2 = {5'd0, _zz_selectReadFifo_0_3};
  assign _zz_selectReadFifo_0_5 = 1'b1;
  assign _zz_selectReadFifo_0_4 = {5'd0, _zz_selectReadFifo_0_5};
  assign _zz_when_ArraySlice_l384 = (_zz_when_ArraySlice_l384_1 % aReg);
  assign _zz_when_ArraySlice_l384_1 = (handshakeTimes_0_value + _zz_when_ArraySlice_l384_2);
  assign _zz_when_ArraySlice_l384_3 = 1'b1;
  assign _zz_when_ArraySlice_l384_2 = {12'd0, _zz_when_ArraySlice_l384_3};
  assign _zz_when_ArraySlice_l389_1 = (selectReadFifo_0 + _zz_when_ArraySlice_l389_2);
  assign _zz_when_ArraySlice_l389_3 = 3'b000;
  assign _zz_when_ArraySlice_l389_2 = {3'd0, _zz_when_ArraySlice_l389_3};
  assign _zz_when_ArraySlice_l389_5 = 1'b1;
  assign _zz_when_ArraySlice_l389_4 = {6'd0, _zz_when_ArraySlice_l389_5};
  assign _zz_when_ArraySlice_l390_1 = (_zz_when_ArraySlice_l390_2 - _zz_when_ArraySlice_l390_3);
  assign _zz_when_ArraySlice_l390 = {7'd0, _zz_when_ArraySlice_l390_1};
  assign _zz_when_ArraySlice_l390_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l390_4 = 1'b1;
  assign _zz_when_ArraySlice_l390_3 = {5'd0, _zz_when_ArraySlice_l390_4};
  assign _zz__zz_when_ArraySlice_l94 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95 = (_zz_when_ArraySlice_l95_1 - _zz_when_ArraySlice_l95_4);
  assign _zz_when_ArraySlice_l95_1 = (_zz_when_ArraySlice_l95_2 + _zz_when_ArraySlice_l95_3);
  assign _zz_when_ArraySlice_l95_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_4 = {1'd0, _zz_when_ArraySlice_l94};
  assign _zz__zz_when_ArraySlice_l392 = (_zz__zz_when_ArraySlice_l392_1 + _zz__zz_when_ArraySlice_l392_2);
  assign _zz__zz_when_ArraySlice_l392_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l392_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l392_3 = {1'd0, _zz_when_ArraySlice_l94};
  assign _zz_when_ArraySlice_l99_1 = 7'h40;
  assign _zz_when_ArraySlice_l99 = _zz_when_ArraySlice_l99_1[5:0];
  assign _zz_when_ArraySlice_l392_8 = (outSliceNumb_0_value + _zz_when_ArraySlice_l392_9);
  assign _zz_when_ArraySlice_l392_10 = 1'b1;
  assign _zz_when_ArraySlice_l392_9 = {6'd0, _zz_when_ArraySlice_l392_10};
  assign _zz_when_ArraySlice_l392_11 = (_zz_when_ArraySlice_l392 / aReg);
  assign _zz_selectReadFifo_0_6 = (selectReadFifo_0 - _zz_selectReadFifo_0_7);
  assign _zz_selectReadFifo_0_7 = {3'd0, bReg};
  assign _zz_selectReadFifo_0_9 = 1'b1;
  assign _zz_selectReadFifo_0_8 = {5'd0, _zz_selectReadFifo_0_9};
  assign _zz_selectReadFifo_0_10 = (selectReadFifo_0 + _zz_selectReadFifo_0_11);
  assign _zz_selectReadFifo_0_11 = (3'b111 * bReg);
  assign _zz_selectReadFifo_0_13 = 1'b1;
  assign _zz_selectReadFifo_0_12 = {5'd0, _zz_selectReadFifo_0_13};
  assign _zz_when_ArraySlice_l165_8 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_8_1);
  assign _zz_when_ArraySlice_l165_8_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_8_1 = {3'd0, _zz_when_ArraySlice_l165_8_2};
  assign _zz_when_ArraySlice_l166_8 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_8_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_8_3);
  assign _zz_when_ArraySlice_l166_8_1 = {1'd0, _zz_when_ArraySlice_l166_8_2};
  assign _zz_when_ArraySlice_l166_8_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_8_4);
  assign _zz_when_ArraySlice_l166_8_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_8_4 = {3'd0, _zz_when_ArraySlice_l166_8_5};
  assign _zz__zz_when_ArraySlice_l112_8 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_8 = (_zz_when_ArraySlice_l113_8_1 - _zz_when_ArraySlice_l113_8_4);
  assign _zz_when_ArraySlice_l113_8_1 = (_zz_when_ArraySlice_l113_8_2 + _zz_when_ArraySlice_l113_8_3);
  assign _zz_when_ArraySlice_l113_8_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_8_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_8_4 = {1'd0, _zz_when_ArraySlice_l112_8};
  assign _zz__zz_when_ArraySlice_l173_8 = (_zz__zz_when_ArraySlice_l173_8_1 + _zz__zz_when_ArraySlice_l173_8_2);
  assign _zz__zz_when_ArraySlice_l173_8_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_8_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_8_3 = {1'd0, _zz_when_ArraySlice_l112_8};
  assign _zz_when_ArraySlice_l118_8_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_8 = _zz_when_ArraySlice_l118_8_1[5:0];
  assign _zz_when_ArraySlice_l173_8_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_8_2 = (_zz_when_ArraySlice_l173_8_3 + _zz_when_ArraySlice_l173_8_8);
  assign _zz_when_ArraySlice_l173_8_3 = (_zz_when_ArraySlice_l173_8 - _zz_when_ArraySlice_l173_8_4);
  assign _zz_when_ArraySlice_l173_8_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_8_6);
  assign _zz_when_ArraySlice_l173_8_4 = {1'd0, _zz_when_ArraySlice_l173_8_5};
  assign _zz_when_ArraySlice_l173_8_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_8_6 = {3'd0, _zz_when_ArraySlice_l173_8_7};
  assign _zz_when_ArraySlice_l173_8_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_9 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_9_1);
  assign _zz_when_ArraySlice_l165_9_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_9_1 = {2'd0, _zz_when_ArraySlice_l165_9_2};
  assign _zz_when_ArraySlice_l166_9 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_9_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_9_2);
  assign _zz_when_ArraySlice_l166_9_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_9_3);
  assign _zz_when_ArraySlice_l166_9_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_9_3 = {2'd0, _zz_when_ArraySlice_l166_9_4};
  assign _zz__zz_when_ArraySlice_l112_9 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_9 = (_zz_when_ArraySlice_l113_9_1 - _zz_when_ArraySlice_l113_9_4);
  assign _zz_when_ArraySlice_l113_9_1 = (_zz_when_ArraySlice_l113_9_2 + _zz_when_ArraySlice_l113_9_3);
  assign _zz_when_ArraySlice_l113_9_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_9_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_9_4 = {1'd0, _zz_when_ArraySlice_l112_9};
  assign _zz__zz_when_ArraySlice_l173_9 = (_zz__zz_when_ArraySlice_l173_9_1 + _zz__zz_when_ArraySlice_l173_9_2);
  assign _zz__zz_when_ArraySlice_l173_9_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_9_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_9_3 = {1'd0, _zz_when_ArraySlice_l112_9};
  assign _zz_when_ArraySlice_l118_9_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_9 = _zz_when_ArraySlice_l118_9_1[5:0];
  assign _zz_when_ArraySlice_l173_9_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_9_1 = {1'd0, _zz_when_ArraySlice_l173_9_2};
  assign _zz_when_ArraySlice_l173_9_3 = (_zz_when_ArraySlice_l173_9_4 + _zz_when_ArraySlice_l173_9_9);
  assign _zz_when_ArraySlice_l173_9_4 = (_zz_when_ArraySlice_l173_9 - _zz_when_ArraySlice_l173_9_5);
  assign _zz_when_ArraySlice_l173_9_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_9_7);
  assign _zz_when_ArraySlice_l173_9_5 = {1'd0, _zz_when_ArraySlice_l173_9_6};
  assign _zz_when_ArraySlice_l173_9_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_9_7 = {2'd0, _zz_when_ArraySlice_l173_9_8};
  assign _zz_when_ArraySlice_l173_9_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_10 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_10_1);
  assign _zz_when_ArraySlice_l165_10_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_10_1 = {1'd0, _zz_when_ArraySlice_l165_10_2};
  assign _zz_when_ArraySlice_l166_10 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_10_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_10_2);
  assign _zz_when_ArraySlice_l166_10_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_10_3);
  assign _zz_when_ArraySlice_l166_10_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_10_3 = {1'd0, _zz_when_ArraySlice_l166_10_4};
  assign _zz__zz_when_ArraySlice_l112_10 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_10 = (_zz_when_ArraySlice_l113_10_1 - _zz_when_ArraySlice_l113_10_4);
  assign _zz_when_ArraySlice_l113_10_1 = (_zz_when_ArraySlice_l113_10_2 + _zz_when_ArraySlice_l113_10_3);
  assign _zz_when_ArraySlice_l113_10_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_10_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_10_4 = {1'd0, _zz_when_ArraySlice_l112_10};
  assign _zz__zz_when_ArraySlice_l173_10 = (_zz__zz_when_ArraySlice_l173_10_1 + _zz__zz_when_ArraySlice_l173_10_2);
  assign _zz__zz_when_ArraySlice_l173_10_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_10_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_10_3 = {1'd0, _zz_when_ArraySlice_l112_10};
  assign _zz_when_ArraySlice_l118_10_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_10 = _zz_when_ArraySlice_l118_10_1[5:0];
  assign _zz_when_ArraySlice_l173_10_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_10_1 = {1'd0, _zz_when_ArraySlice_l173_10_2};
  assign _zz_when_ArraySlice_l173_10_3 = (_zz_when_ArraySlice_l173_10_4 + _zz_when_ArraySlice_l173_10_9);
  assign _zz_when_ArraySlice_l173_10_4 = (_zz_when_ArraySlice_l173_10 - _zz_when_ArraySlice_l173_10_5);
  assign _zz_when_ArraySlice_l173_10_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_10_7);
  assign _zz_when_ArraySlice_l173_10_5 = {1'd0, _zz_when_ArraySlice_l173_10_6};
  assign _zz_when_ArraySlice_l173_10_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_10_7 = {1'd0, _zz_when_ArraySlice_l173_10_8};
  assign _zz_when_ArraySlice_l173_10_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_11 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_11_1);
  assign _zz_when_ArraySlice_l165_11_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_11_1 = {1'd0, _zz_when_ArraySlice_l165_11_2};
  assign _zz_when_ArraySlice_l166_11 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_11_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_11_2);
  assign _zz_when_ArraySlice_l166_11_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_11_3);
  assign _zz_when_ArraySlice_l166_11_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_11_3 = {1'd0, _zz_when_ArraySlice_l166_11_4};
  assign _zz__zz_when_ArraySlice_l112_11 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_11 = (_zz_when_ArraySlice_l113_11_1 - _zz_when_ArraySlice_l113_11_4);
  assign _zz_when_ArraySlice_l113_11_1 = (_zz_when_ArraySlice_l113_11_2 + _zz_when_ArraySlice_l113_11_3);
  assign _zz_when_ArraySlice_l113_11_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_11_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_11_4 = {1'd0, _zz_when_ArraySlice_l112_11};
  assign _zz__zz_when_ArraySlice_l173_11 = (_zz__zz_when_ArraySlice_l173_11_1 + _zz__zz_when_ArraySlice_l173_11_2);
  assign _zz__zz_when_ArraySlice_l173_11_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_11_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_11_3 = {1'd0, _zz_when_ArraySlice_l112_11};
  assign _zz_when_ArraySlice_l118_11_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_11 = _zz_when_ArraySlice_l118_11_1[5:0];
  assign _zz_when_ArraySlice_l173_11_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_11_1 = {1'd0, _zz_when_ArraySlice_l173_11_2};
  assign _zz_when_ArraySlice_l173_11_3 = (_zz_when_ArraySlice_l173_11_4 + _zz_when_ArraySlice_l173_11_9);
  assign _zz_when_ArraySlice_l173_11_4 = (_zz_when_ArraySlice_l173_11 - _zz_when_ArraySlice_l173_11_5);
  assign _zz_when_ArraySlice_l173_11_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_11_7);
  assign _zz_when_ArraySlice_l173_11_5 = {1'd0, _zz_when_ArraySlice_l173_11_6};
  assign _zz_when_ArraySlice_l173_11_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_11_7 = {1'd0, _zz_when_ArraySlice_l173_11_8};
  assign _zz_when_ArraySlice_l173_11_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_12 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_12_1);
  assign _zz_when_ArraySlice_l165_12_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_12 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_12_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_12_2);
  assign _zz_when_ArraySlice_l166_12_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_12_3);
  assign _zz_when_ArraySlice_l166_12_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_12 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_12 = (_zz_when_ArraySlice_l113_12_1 - _zz_when_ArraySlice_l113_12_4);
  assign _zz_when_ArraySlice_l113_12_1 = (_zz_when_ArraySlice_l113_12_2 + _zz_when_ArraySlice_l113_12_3);
  assign _zz_when_ArraySlice_l113_12_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_12_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_12_4 = {1'd0, _zz_when_ArraySlice_l112_12};
  assign _zz__zz_when_ArraySlice_l173_12 = (_zz__zz_when_ArraySlice_l173_12_1 + _zz__zz_when_ArraySlice_l173_12_2);
  assign _zz__zz_when_ArraySlice_l173_12_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_12_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_12_3 = {1'd0, _zz_when_ArraySlice_l112_12};
  assign _zz_when_ArraySlice_l118_12_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_12 = _zz_when_ArraySlice_l118_12_1[5:0];
  assign _zz_when_ArraySlice_l173_12_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_12_1 = {1'd0, _zz_when_ArraySlice_l173_12_2};
  assign _zz_when_ArraySlice_l173_12_3 = (_zz_when_ArraySlice_l173_12_4 + _zz_when_ArraySlice_l173_12_8);
  assign _zz_when_ArraySlice_l173_12_4 = (_zz_when_ArraySlice_l173_12 - _zz_when_ArraySlice_l173_12_5);
  assign _zz_when_ArraySlice_l173_12_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_12_7);
  assign _zz_when_ArraySlice_l173_12_5 = {1'd0, _zz_when_ArraySlice_l173_12_6};
  assign _zz_when_ArraySlice_l173_12_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_12_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_13 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_13_1);
  assign _zz_when_ArraySlice_l165_13_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_13_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_13 = {1'd0, _zz_when_ArraySlice_l166_13_1};
  assign _zz_when_ArraySlice_l166_13_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_13_3);
  assign _zz_when_ArraySlice_l166_13_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_13_4);
  assign _zz_when_ArraySlice_l166_13_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_13 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_13 = (_zz_when_ArraySlice_l113_13_1 - _zz_when_ArraySlice_l113_13_4);
  assign _zz_when_ArraySlice_l113_13_1 = (_zz_when_ArraySlice_l113_13_2 + _zz_when_ArraySlice_l113_13_3);
  assign _zz_when_ArraySlice_l113_13_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_13_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_13_4 = {1'd0, _zz_when_ArraySlice_l112_13};
  assign _zz__zz_when_ArraySlice_l173_13 = (_zz__zz_when_ArraySlice_l173_13_1 + _zz__zz_when_ArraySlice_l173_13_2);
  assign _zz__zz_when_ArraySlice_l173_13_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_13_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_13_3 = {1'd0, _zz_when_ArraySlice_l112_13};
  assign _zz_when_ArraySlice_l118_13_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_13 = _zz_when_ArraySlice_l118_13_1[5:0];
  assign _zz_when_ArraySlice_l173_13_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_13_1 = {2'd0, _zz_when_ArraySlice_l173_13_2};
  assign _zz_when_ArraySlice_l173_13_3 = (_zz_when_ArraySlice_l173_13_4 + _zz_when_ArraySlice_l173_13_8);
  assign _zz_when_ArraySlice_l173_13_4 = (_zz_when_ArraySlice_l173_13 - _zz_when_ArraySlice_l173_13_5);
  assign _zz_when_ArraySlice_l173_13_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_13_7);
  assign _zz_when_ArraySlice_l173_13_5 = {1'd0, _zz_when_ArraySlice_l173_13_6};
  assign _zz_when_ArraySlice_l173_13_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_13_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_14 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_14_1);
  assign _zz_when_ArraySlice_l165_14_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_14_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_14 = {1'd0, _zz_when_ArraySlice_l166_14_1};
  assign _zz_when_ArraySlice_l166_14_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_14_3);
  assign _zz_when_ArraySlice_l166_14_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_14_4);
  assign _zz_when_ArraySlice_l166_14_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_14 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_14 = (_zz_when_ArraySlice_l113_14_1 - _zz_when_ArraySlice_l113_14_4);
  assign _zz_when_ArraySlice_l113_14_1 = (_zz_when_ArraySlice_l113_14_2 + _zz_when_ArraySlice_l113_14_3);
  assign _zz_when_ArraySlice_l113_14_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_14_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_14_4 = {1'd0, _zz_when_ArraySlice_l112_14};
  assign _zz__zz_when_ArraySlice_l173_14 = (_zz__zz_when_ArraySlice_l173_14_1 + _zz__zz_when_ArraySlice_l173_14_2);
  assign _zz__zz_when_ArraySlice_l173_14_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_14_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_14_3 = {1'd0, _zz_when_ArraySlice_l112_14};
  assign _zz_when_ArraySlice_l118_14_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_14 = _zz_when_ArraySlice_l118_14_1[5:0];
  assign _zz_when_ArraySlice_l173_14_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_14_1 = {2'd0, _zz_when_ArraySlice_l173_14_2};
  assign _zz_when_ArraySlice_l173_14_3 = (_zz_when_ArraySlice_l173_14_4 + _zz_when_ArraySlice_l173_14_8);
  assign _zz_when_ArraySlice_l173_14_4 = (_zz_when_ArraySlice_l173_14 - _zz_when_ArraySlice_l173_14_5);
  assign _zz_when_ArraySlice_l173_14_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_14_7);
  assign _zz_when_ArraySlice_l173_14_5 = {1'd0, _zz_when_ArraySlice_l173_14_6};
  assign _zz_when_ArraySlice_l173_14_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_14_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_15 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_15_1);
  assign _zz_when_ArraySlice_l165_15_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_15_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_15 = {2'd0, _zz_when_ArraySlice_l166_15_1};
  assign _zz_when_ArraySlice_l166_15_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_15_3);
  assign _zz_when_ArraySlice_l166_15_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_15_4);
  assign _zz_when_ArraySlice_l166_15_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_15 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_15 = (_zz_when_ArraySlice_l113_15_1 - _zz_when_ArraySlice_l113_15_4);
  assign _zz_when_ArraySlice_l113_15_1 = (_zz_when_ArraySlice_l113_15_2 + _zz_when_ArraySlice_l113_15_3);
  assign _zz_when_ArraySlice_l113_15_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_15_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_15_4 = {1'd0, _zz_when_ArraySlice_l112_15};
  assign _zz__zz_when_ArraySlice_l173_15 = (_zz__zz_when_ArraySlice_l173_15_1 + _zz__zz_when_ArraySlice_l173_15_2);
  assign _zz__zz_when_ArraySlice_l173_15_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_15_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_15_3 = {1'd0, _zz_when_ArraySlice_l112_15};
  assign _zz_when_ArraySlice_l118_15_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_15 = _zz_when_ArraySlice_l118_15_1[5:0];
  assign _zz_when_ArraySlice_l173_15_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_15_1 = {3'd0, _zz_when_ArraySlice_l173_15_2};
  assign _zz_when_ArraySlice_l173_15_3 = (_zz_when_ArraySlice_l173_15_4 + _zz_when_ArraySlice_l173_15_8);
  assign _zz_when_ArraySlice_l173_15_4 = (_zz_when_ArraySlice_l173_15 - _zz_when_ArraySlice_l173_15_5);
  assign _zz_when_ArraySlice_l173_15_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_15_7);
  assign _zz_when_ArraySlice_l173_15_5 = {1'd0, _zz_when_ArraySlice_l173_15_6};
  assign _zz_when_ArraySlice_l173_15_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_15_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l401 = (_zz_when_ArraySlice_l401_1 + _zz_when_ArraySlice_l401_6);
  assign _zz_when_ArraySlice_l401_1 = (_zz_when_ArraySlice_l401_2 + _zz_when_ArraySlice_l401_4);
  assign _zz_when_ArraySlice_l401_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l401_3);
  assign _zz_when_ArraySlice_l401_3 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l401_5 = 1'b1;
  assign _zz_when_ArraySlice_l401_4 = {5'd0, _zz_when_ArraySlice_l401_5};
  assign _zz_when_ArraySlice_l401_7 = 3'b000;
  assign _zz_when_ArraySlice_l401_6 = {3'd0, _zz_when_ArraySlice_l401_7};
  assign _zz_selectReadFifo_0_15 = 1'b1;
  assign _zz_selectReadFifo_0_14 = {5'd0, _zz_selectReadFifo_0_15};
  assign _zz_when_ArraySlice_l405 = (_zz_when_ArraySlice_l405_1 % aReg);
  assign _zz_when_ArraySlice_l405_1 = (handshakeTimes_0_value + _zz_when_ArraySlice_l405_2);
  assign _zz_when_ArraySlice_l405_3 = 1'b1;
  assign _zz_when_ArraySlice_l405_2 = {12'd0, _zz_when_ArraySlice_l405_3};
  assign _zz_when_ArraySlice_l409_1 = (selectReadFifo_0 + _zz_when_ArraySlice_l409_2);
  assign _zz_when_ArraySlice_l409_3 = 3'b000;
  assign _zz_when_ArraySlice_l409_2 = {3'd0, _zz_when_ArraySlice_l409_3};
  assign _zz_when_ArraySlice_l410_1 = (_zz_when_ArraySlice_l410_2 - _zz_when_ArraySlice_l410_3);
  assign _zz_when_ArraySlice_l410 = {7'd0, _zz_when_ArraySlice_l410_1};
  assign _zz_when_ArraySlice_l410_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l410_4 = 1'b1;
  assign _zz_when_ArraySlice_l410_3 = {5'd0, _zz_when_ArraySlice_l410_4};
  assign _zz__zz_when_ArraySlice_l94_1 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_1_1 = (_zz_when_ArraySlice_l95_1_2 - _zz_when_ArraySlice_l95_1_5);
  assign _zz_when_ArraySlice_l95_1_2 = (_zz_when_ArraySlice_l95_1_3 + _zz_when_ArraySlice_l95_1_4);
  assign _zz_when_ArraySlice_l95_1_3 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_1_4 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_1_5 = {1'd0, _zz_when_ArraySlice_l94_1};
  assign _zz__zz_when_ArraySlice_l412 = (_zz__zz_when_ArraySlice_l412_1 + _zz__zz_when_ArraySlice_l412_2);
  assign _zz__zz_when_ArraySlice_l412_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l412_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l412_3 = {1'd0, _zz_when_ArraySlice_l94_1};
  assign _zz_when_ArraySlice_l99_1_2 = 7'h40;
  assign _zz_when_ArraySlice_l99_1_1 = _zz_when_ArraySlice_l99_1_2[5:0];
  assign _zz_when_ArraySlice_l412_8 = (outSliceNumb_0_value + _zz_when_ArraySlice_l412_9);
  assign _zz_when_ArraySlice_l412_10 = 1'b1;
  assign _zz_when_ArraySlice_l412_9 = {6'd0, _zz_when_ArraySlice_l412_10};
  assign _zz_when_ArraySlice_l412_11 = (_zz_when_ArraySlice_l412 / aReg);
  assign _zz_selectReadFifo_0_16 = (selectReadFifo_0 - _zz_selectReadFifo_0_17);
  assign _zz_selectReadFifo_0_17 = {3'd0, bReg};
  assign _zz_selectReadFifo_0_19 = 1'b1;
  assign _zz_selectReadFifo_0_18 = {5'd0, _zz_selectReadFifo_0_19};
  assign _zz_selectReadFifo_0_20 = (selectReadFifo_0 + _zz_selectReadFifo_0_21);
  assign _zz_selectReadFifo_0_21 = (3'b111 * bReg);
  assign _zz_selectReadFifo_0_23 = 1'b1;
  assign _zz_selectReadFifo_0_22 = {5'd0, _zz_selectReadFifo_0_23};
  assign _zz_when_ArraySlice_l165_16 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_16_1);
  assign _zz_when_ArraySlice_l165_16_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_16_1 = {3'd0, _zz_when_ArraySlice_l165_16_2};
  assign _zz_when_ArraySlice_l166_16 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_16_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_16_3);
  assign _zz_when_ArraySlice_l166_16_1 = {1'd0, _zz_when_ArraySlice_l166_16_2};
  assign _zz_when_ArraySlice_l166_16_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_16_4);
  assign _zz_when_ArraySlice_l166_16_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_16_4 = {3'd0, _zz_when_ArraySlice_l166_16_5};
  assign _zz__zz_when_ArraySlice_l112_16 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_16 = (_zz_when_ArraySlice_l113_16_1 - _zz_when_ArraySlice_l113_16_4);
  assign _zz_when_ArraySlice_l113_16_1 = (_zz_when_ArraySlice_l113_16_2 + _zz_when_ArraySlice_l113_16_3);
  assign _zz_when_ArraySlice_l113_16_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_16_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_16_4 = {1'd0, _zz_when_ArraySlice_l112_16};
  assign _zz__zz_when_ArraySlice_l173_16 = (_zz__zz_when_ArraySlice_l173_16_1 + _zz__zz_when_ArraySlice_l173_16_2);
  assign _zz__zz_when_ArraySlice_l173_16_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_16_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_16_3 = {1'd0, _zz_when_ArraySlice_l112_16};
  assign _zz_when_ArraySlice_l118_16_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_16 = _zz_when_ArraySlice_l118_16_1[5:0];
  assign _zz_when_ArraySlice_l173_16_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_16_2 = (_zz_when_ArraySlice_l173_16_3 + _zz_when_ArraySlice_l173_16_8);
  assign _zz_when_ArraySlice_l173_16_3 = (_zz_when_ArraySlice_l173_16 - _zz_when_ArraySlice_l173_16_4);
  assign _zz_when_ArraySlice_l173_16_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_16_6);
  assign _zz_when_ArraySlice_l173_16_4 = {1'd0, _zz_when_ArraySlice_l173_16_5};
  assign _zz_when_ArraySlice_l173_16_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_16_6 = {3'd0, _zz_when_ArraySlice_l173_16_7};
  assign _zz_when_ArraySlice_l173_16_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_17 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_17_1);
  assign _zz_when_ArraySlice_l165_17_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_17_1 = {2'd0, _zz_when_ArraySlice_l165_17_2};
  assign _zz_when_ArraySlice_l166_17 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_17_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_17_2);
  assign _zz_when_ArraySlice_l166_17_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_17_3);
  assign _zz_when_ArraySlice_l166_17_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_17_3 = {2'd0, _zz_when_ArraySlice_l166_17_4};
  assign _zz__zz_when_ArraySlice_l112_17 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_17 = (_zz_when_ArraySlice_l113_17_1 - _zz_when_ArraySlice_l113_17_4);
  assign _zz_when_ArraySlice_l113_17_1 = (_zz_when_ArraySlice_l113_17_2 + _zz_when_ArraySlice_l113_17_3);
  assign _zz_when_ArraySlice_l113_17_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_17_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_17_4 = {1'd0, _zz_when_ArraySlice_l112_17};
  assign _zz__zz_when_ArraySlice_l173_17 = (_zz__zz_when_ArraySlice_l173_17_1 + _zz__zz_when_ArraySlice_l173_17_2);
  assign _zz__zz_when_ArraySlice_l173_17_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_17_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_17_3 = {1'd0, _zz_when_ArraySlice_l112_17};
  assign _zz_when_ArraySlice_l118_17_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_17 = _zz_when_ArraySlice_l118_17_1[5:0];
  assign _zz_when_ArraySlice_l173_17_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_17_1 = {1'd0, _zz_when_ArraySlice_l173_17_2};
  assign _zz_when_ArraySlice_l173_17_3 = (_zz_when_ArraySlice_l173_17_4 + _zz_when_ArraySlice_l173_17_9);
  assign _zz_when_ArraySlice_l173_17_4 = (_zz_when_ArraySlice_l173_17 - _zz_when_ArraySlice_l173_17_5);
  assign _zz_when_ArraySlice_l173_17_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_17_7);
  assign _zz_when_ArraySlice_l173_17_5 = {1'd0, _zz_when_ArraySlice_l173_17_6};
  assign _zz_when_ArraySlice_l173_17_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_17_7 = {2'd0, _zz_when_ArraySlice_l173_17_8};
  assign _zz_when_ArraySlice_l173_17_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_18 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_18_1);
  assign _zz_when_ArraySlice_l165_18_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_18_1 = {1'd0, _zz_when_ArraySlice_l165_18_2};
  assign _zz_when_ArraySlice_l166_18 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_18_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_18_2);
  assign _zz_when_ArraySlice_l166_18_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_18_3);
  assign _zz_when_ArraySlice_l166_18_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_18_3 = {1'd0, _zz_when_ArraySlice_l166_18_4};
  assign _zz__zz_when_ArraySlice_l112_18 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_18 = (_zz_when_ArraySlice_l113_18_1 - _zz_when_ArraySlice_l113_18_4);
  assign _zz_when_ArraySlice_l113_18_1 = (_zz_when_ArraySlice_l113_18_2 + _zz_when_ArraySlice_l113_18_3);
  assign _zz_when_ArraySlice_l113_18_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_18_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_18_4 = {1'd0, _zz_when_ArraySlice_l112_18};
  assign _zz__zz_when_ArraySlice_l173_18 = (_zz__zz_when_ArraySlice_l173_18_1 + _zz__zz_when_ArraySlice_l173_18_2);
  assign _zz__zz_when_ArraySlice_l173_18_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_18_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_18_3 = {1'd0, _zz_when_ArraySlice_l112_18};
  assign _zz_when_ArraySlice_l118_18_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_18 = _zz_when_ArraySlice_l118_18_1[5:0];
  assign _zz_when_ArraySlice_l173_18_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_18_1 = {1'd0, _zz_when_ArraySlice_l173_18_2};
  assign _zz_when_ArraySlice_l173_18_3 = (_zz_when_ArraySlice_l173_18_4 + _zz_when_ArraySlice_l173_18_9);
  assign _zz_when_ArraySlice_l173_18_4 = (_zz_when_ArraySlice_l173_18 - _zz_when_ArraySlice_l173_18_5);
  assign _zz_when_ArraySlice_l173_18_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_18_7);
  assign _zz_when_ArraySlice_l173_18_5 = {1'd0, _zz_when_ArraySlice_l173_18_6};
  assign _zz_when_ArraySlice_l173_18_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_18_7 = {1'd0, _zz_when_ArraySlice_l173_18_8};
  assign _zz_when_ArraySlice_l173_18_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_19 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_19_1);
  assign _zz_when_ArraySlice_l165_19_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_19_1 = {1'd0, _zz_when_ArraySlice_l165_19_2};
  assign _zz_when_ArraySlice_l166_19 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_19_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_19_2);
  assign _zz_when_ArraySlice_l166_19_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_19_3);
  assign _zz_when_ArraySlice_l166_19_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_19_3 = {1'd0, _zz_when_ArraySlice_l166_19_4};
  assign _zz__zz_when_ArraySlice_l112_19 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_19 = (_zz_when_ArraySlice_l113_19_1 - _zz_when_ArraySlice_l113_19_4);
  assign _zz_when_ArraySlice_l113_19_1 = (_zz_when_ArraySlice_l113_19_2 + _zz_when_ArraySlice_l113_19_3);
  assign _zz_when_ArraySlice_l113_19_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_19_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_19_4 = {1'd0, _zz_when_ArraySlice_l112_19};
  assign _zz__zz_when_ArraySlice_l173_19 = (_zz__zz_when_ArraySlice_l173_19_1 + _zz__zz_when_ArraySlice_l173_19_2);
  assign _zz__zz_when_ArraySlice_l173_19_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_19_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_19_3 = {1'd0, _zz_when_ArraySlice_l112_19};
  assign _zz_when_ArraySlice_l118_19_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_19 = _zz_when_ArraySlice_l118_19_1[5:0];
  assign _zz_when_ArraySlice_l173_19_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_19_1 = {1'd0, _zz_when_ArraySlice_l173_19_2};
  assign _zz_when_ArraySlice_l173_19_3 = (_zz_when_ArraySlice_l173_19_4 + _zz_when_ArraySlice_l173_19_9);
  assign _zz_when_ArraySlice_l173_19_4 = (_zz_when_ArraySlice_l173_19 - _zz_when_ArraySlice_l173_19_5);
  assign _zz_when_ArraySlice_l173_19_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_19_7);
  assign _zz_when_ArraySlice_l173_19_5 = {1'd0, _zz_when_ArraySlice_l173_19_6};
  assign _zz_when_ArraySlice_l173_19_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_19_7 = {1'd0, _zz_when_ArraySlice_l173_19_8};
  assign _zz_when_ArraySlice_l173_19_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_20 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_20_1);
  assign _zz_when_ArraySlice_l165_20_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_20 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_20_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_20_2);
  assign _zz_when_ArraySlice_l166_20_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_20_3);
  assign _zz_when_ArraySlice_l166_20_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_20 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_20 = (_zz_when_ArraySlice_l113_20_1 - _zz_when_ArraySlice_l113_20_4);
  assign _zz_when_ArraySlice_l113_20_1 = (_zz_when_ArraySlice_l113_20_2 + _zz_when_ArraySlice_l113_20_3);
  assign _zz_when_ArraySlice_l113_20_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_20_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_20_4 = {1'd0, _zz_when_ArraySlice_l112_20};
  assign _zz__zz_when_ArraySlice_l173_20 = (_zz__zz_when_ArraySlice_l173_20_1 + _zz__zz_when_ArraySlice_l173_20_2);
  assign _zz__zz_when_ArraySlice_l173_20_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_20_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_20_3 = {1'd0, _zz_when_ArraySlice_l112_20};
  assign _zz_when_ArraySlice_l118_20_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_20 = _zz_when_ArraySlice_l118_20_1[5:0];
  assign _zz_when_ArraySlice_l173_20_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_20_1 = {1'd0, _zz_when_ArraySlice_l173_20_2};
  assign _zz_when_ArraySlice_l173_20_3 = (_zz_when_ArraySlice_l173_20_4 + _zz_when_ArraySlice_l173_20_8);
  assign _zz_when_ArraySlice_l173_20_4 = (_zz_when_ArraySlice_l173_20 - _zz_when_ArraySlice_l173_20_5);
  assign _zz_when_ArraySlice_l173_20_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_20_7);
  assign _zz_when_ArraySlice_l173_20_5 = {1'd0, _zz_when_ArraySlice_l173_20_6};
  assign _zz_when_ArraySlice_l173_20_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_20_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_21 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_21_1);
  assign _zz_when_ArraySlice_l165_21_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_21_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_21 = {1'd0, _zz_when_ArraySlice_l166_21_1};
  assign _zz_when_ArraySlice_l166_21_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_21_3);
  assign _zz_when_ArraySlice_l166_21_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_21_4);
  assign _zz_when_ArraySlice_l166_21_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_21 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_21 = (_zz_when_ArraySlice_l113_21_1 - _zz_when_ArraySlice_l113_21_4);
  assign _zz_when_ArraySlice_l113_21_1 = (_zz_when_ArraySlice_l113_21_2 + _zz_when_ArraySlice_l113_21_3);
  assign _zz_when_ArraySlice_l113_21_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_21_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_21_4 = {1'd0, _zz_when_ArraySlice_l112_21};
  assign _zz__zz_when_ArraySlice_l173_21 = (_zz__zz_when_ArraySlice_l173_21_1 + _zz__zz_when_ArraySlice_l173_21_2);
  assign _zz__zz_when_ArraySlice_l173_21_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_21_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_21_3 = {1'd0, _zz_when_ArraySlice_l112_21};
  assign _zz_when_ArraySlice_l118_21_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_21 = _zz_when_ArraySlice_l118_21_1[5:0];
  assign _zz_when_ArraySlice_l173_21_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_21_1 = {2'd0, _zz_when_ArraySlice_l173_21_2};
  assign _zz_when_ArraySlice_l173_21_3 = (_zz_when_ArraySlice_l173_21_4 + _zz_when_ArraySlice_l173_21_8);
  assign _zz_when_ArraySlice_l173_21_4 = (_zz_when_ArraySlice_l173_21 - _zz_when_ArraySlice_l173_21_5);
  assign _zz_when_ArraySlice_l173_21_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_21_7);
  assign _zz_when_ArraySlice_l173_21_5 = {1'd0, _zz_when_ArraySlice_l173_21_6};
  assign _zz_when_ArraySlice_l173_21_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_21_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_22 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_22_1);
  assign _zz_when_ArraySlice_l165_22_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_22_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_22 = {1'd0, _zz_when_ArraySlice_l166_22_1};
  assign _zz_when_ArraySlice_l166_22_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_22_3);
  assign _zz_when_ArraySlice_l166_22_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_22_4);
  assign _zz_when_ArraySlice_l166_22_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_22 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_22 = (_zz_when_ArraySlice_l113_22_1 - _zz_when_ArraySlice_l113_22_4);
  assign _zz_when_ArraySlice_l113_22_1 = (_zz_when_ArraySlice_l113_22_2 + _zz_when_ArraySlice_l113_22_3);
  assign _zz_when_ArraySlice_l113_22_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_22_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_22_4 = {1'd0, _zz_when_ArraySlice_l112_22};
  assign _zz__zz_when_ArraySlice_l173_22 = (_zz__zz_when_ArraySlice_l173_22_1 + _zz__zz_when_ArraySlice_l173_22_2);
  assign _zz__zz_when_ArraySlice_l173_22_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_22_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_22_3 = {1'd0, _zz_when_ArraySlice_l112_22};
  assign _zz_when_ArraySlice_l118_22_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_22 = _zz_when_ArraySlice_l118_22_1[5:0];
  assign _zz_when_ArraySlice_l173_22_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_22_1 = {2'd0, _zz_when_ArraySlice_l173_22_2};
  assign _zz_when_ArraySlice_l173_22_3 = (_zz_when_ArraySlice_l173_22_4 + _zz_when_ArraySlice_l173_22_8);
  assign _zz_when_ArraySlice_l173_22_4 = (_zz_when_ArraySlice_l173_22 - _zz_when_ArraySlice_l173_22_5);
  assign _zz_when_ArraySlice_l173_22_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_22_7);
  assign _zz_when_ArraySlice_l173_22_5 = {1'd0, _zz_when_ArraySlice_l173_22_6};
  assign _zz_when_ArraySlice_l173_22_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_22_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_23 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_23_1);
  assign _zz_when_ArraySlice_l165_23_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_23_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_23 = {2'd0, _zz_when_ArraySlice_l166_23_1};
  assign _zz_when_ArraySlice_l166_23_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_23_3);
  assign _zz_when_ArraySlice_l166_23_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_23_4);
  assign _zz_when_ArraySlice_l166_23_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_23 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_23 = (_zz_when_ArraySlice_l113_23_1 - _zz_when_ArraySlice_l113_23_4);
  assign _zz_when_ArraySlice_l113_23_1 = (_zz_when_ArraySlice_l113_23_2 + _zz_when_ArraySlice_l113_23_3);
  assign _zz_when_ArraySlice_l113_23_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_23_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_23_4 = {1'd0, _zz_when_ArraySlice_l112_23};
  assign _zz__zz_when_ArraySlice_l173_23 = (_zz__zz_when_ArraySlice_l173_23_1 + _zz__zz_when_ArraySlice_l173_23_2);
  assign _zz__zz_when_ArraySlice_l173_23_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_23_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_23_3 = {1'd0, _zz_when_ArraySlice_l112_23};
  assign _zz_when_ArraySlice_l118_23_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_23 = _zz_when_ArraySlice_l118_23_1[5:0];
  assign _zz_when_ArraySlice_l173_23_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_23_1 = {3'd0, _zz_when_ArraySlice_l173_23_2};
  assign _zz_when_ArraySlice_l173_23_3 = (_zz_when_ArraySlice_l173_23_4 + _zz_when_ArraySlice_l173_23_8);
  assign _zz_when_ArraySlice_l173_23_4 = (_zz_when_ArraySlice_l173_23 - _zz_when_ArraySlice_l173_23_5);
  assign _zz_when_ArraySlice_l173_23_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_23_7);
  assign _zz_when_ArraySlice_l173_23_5 = {1'd0, _zz_when_ArraySlice_l173_23_6};
  assign _zz_when_ArraySlice_l173_23_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_23_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l421 = (_zz_when_ArraySlice_l421_1 + _zz_when_ArraySlice_l421_6);
  assign _zz_when_ArraySlice_l421_1 = (_zz_when_ArraySlice_l421_2 + _zz_when_ArraySlice_l421_4);
  assign _zz_when_ArraySlice_l421_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l421_3);
  assign _zz_when_ArraySlice_l421_3 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l421_5 = 1'b1;
  assign _zz_when_ArraySlice_l421_4 = {5'd0, _zz_when_ArraySlice_l421_5};
  assign _zz_when_ArraySlice_l421_7 = 3'b000;
  assign _zz_when_ArraySlice_l421_6 = {3'd0, _zz_when_ArraySlice_l421_7};
  assign _zz_selectReadFifo_0_25 = 1'b1;
  assign _zz_selectReadFifo_0_24 = {5'd0, _zz_selectReadFifo_0_25};
  assign _zz_when_ArraySlice_l425 = (_zz_when_ArraySlice_l425_1 % aReg);
  assign _zz_when_ArraySlice_l425_1 = (handshakeTimes_0_value + _zz_when_ArraySlice_l425_2);
  assign _zz_when_ArraySlice_l425_3 = 1'b1;
  assign _zz_when_ArraySlice_l425_2 = {12'd0, _zz_when_ArraySlice_l425_3};
  assign _zz_when_ArraySlice_l436_1 = (_zz_when_ArraySlice_l436_2 - _zz_when_ArraySlice_l436_3);
  assign _zz_when_ArraySlice_l436 = {7'd0, _zz_when_ArraySlice_l436_1};
  assign _zz_when_ArraySlice_l436_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l436_4 = 1'b1;
  assign _zz_when_ArraySlice_l436_3 = {5'd0, _zz_when_ArraySlice_l436_4};
  assign _zz__zz_when_ArraySlice_l94_2 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_2_1 = (_zz_when_ArraySlice_l95_2_2 - _zz_when_ArraySlice_l95_2_5);
  assign _zz_when_ArraySlice_l95_2_2 = (_zz_when_ArraySlice_l95_2_3 + _zz_when_ArraySlice_l95_2_4);
  assign _zz_when_ArraySlice_l95_2_3 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_2_4 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_2_5 = {1'd0, _zz_when_ArraySlice_l94_2};
  assign _zz__zz_when_ArraySlice_l437 = (_zz__zz_when_ArraySlice_l437_1 + _zz__zz_when_ArraySlice_l437_2);
  assign _zz__zz_when_ArraySlice_l437_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l437_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l437_3 = {1'd0, _zz_when_ArraySlice_l94_2};
  assign _zz_when_ArraySlice_l99_2_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_2 = _zz_when_ArraySlice_l99_2_1[5:0];
  assign _zz_when_ArraySlice_l437_8 = (outSliceNumb_0_value + _zz_when_ArraySlice_l437_9);
  assign _zz_when_ArraySlice_l437_10 = 1'b1;
  assign _zz_when_ArraySlice_l437_9 = {6'd0, _zz_when_ArraySlice_l437_10};
  assign _zz_when_ArraySlice_l437_11 = (_zz_when_ArraySlice_l437 / aReg);
  assign _zz_selectReadFifo_0_26 = (selectReadFifo_0 - _zz_selectReadFifo_0_27);
  assign _zz_selectReadFifo_0_27 = {3'd0, bReg};
  assign _zz_selectReadFifo_0_29 = 1'b1;
  assign _zz_selectReadFifo_0_28 = {5'd0, _zz_selectReadFifo_0_29};
  assign _zz_when_ArraySlice_l165_24 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_24_1);
  assign _zz_when_ArraySlice_l165_24_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_24_1 = {3'd0, _zz_when_ArraySlice_l165_24_2};
  assign _zz_when_ArraySlice_l166_24 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_24_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_24_3);
  assign _zz_when_ArraySlice_l166_24_1 = {1'd0, _zz_when_ArraySlice_l166_24_2};
  assign _zz_when_ArraySlice_l166_24_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_24_4);
  assign _zz_when_ArraySlice_l166_24_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_24_4 = {3'd0, _zz_when_ArraySlice_l166_24_5};
  assign _zz__zz_when_ArraySlice_l112_24 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_24 = (_zz_when_ArraySlice_l113_24_1 - _zz_when_ArraySlice_l113_24_4);
  assign _zz_when_ArraySlice_l113_24_1 = (_zz_when_ArraySlice_l113_24_2 + _zz_when_ArraySlice_l113_24_3);
  assign _zz_when_ArraySlice_l113_24_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_24_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_24_4 = {1'd0, _zz_when_ArraySlice_l112_24};
  assign _zz__zz_when_ArraySlice_l173_24 = (_zz__zz_when_ArraySlice_l173_24_1 + _zz__zz_when_ArraySlice_l173_24_2);
  assign _zz__zz_when_ArraySlice_l173_24_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_24_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_24_3 = {1'd0, _zz_when_ArraySlice_l112_24};
  assign _zz_when_ArraySlice_l118_24_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_24 = _zz_when_ArraySlice_l118_24_1[5:0];
  assign _zz_when_ArraySlice_l173_24_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_24_2 = (_zz_when_ArraySlice_l173_24_3 + _zz_when_ArraySlice_l173_24_8);
  assign _zz_when_ArraySlice_l173_24_3 = (_zz_when_ArraySlice_l173_24 - _zz_when_ArraySlice_l173_24_4);
  assign _zz_when_ArraySlice_l173_24_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_24_6);
  assign _zz_when_ArraySlice_l173_24_4 = {1'd0, _zz_when_ArraySlice_l173_24_5};
  assign _zz_when_ArraySlice_l173_24_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_24_6 = {3'd0, _zz_when_ArraySlice_l173_24_7};
  assign _zz_when_ArraySlice_l173_24_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_25 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_25_1);
  assign _zz_when_ArraySlice_l165_25_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_25_1 = {2'd0, _zz_when_ArraySlice_l165_25_2};
  assign _zz_when_ArraySlice_l166_25 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_25_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_25_2);
  assign _zz_when_ArraySlice_l166_25_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_25_3);
  assign _zz_when_ArraySlice_l166_25_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_25_3 = {2'd0, _zz_when_ArraySlice_l166_25_4};
  assign _zz__zz_when_ArraySlice_l112_25 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_25 = (_zz_when_ArraySlice_l113_25_1 - _zz_when_ArraySlice_l113_25_4);
  assign _zz_when_ArraySlice_l113_25_1 = (_zz_when_ArraySlice_l113_25_2 + _zz_when_ArraySlice_l113_25_3);
  assign _zz_when_ArraySlice_l113_25_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_25_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_25_4 = {1'd0, _zz_when_ArraySlice_l112_25};
  assign _zz__zz_when_ArraySlice_l173_25 = (_zz__zz_when_ArraySlice_l173_25_1 + _zz__zz_when_ArraySlice_l173_25_2);
  assign _zz__zz_when_ArraySlice_l173_25_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_25_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_25_3 = {1'd0, _zz_when_ArraySlice_l112_25};
  assign _zz_when_ArraySlice_l118_25_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_25 = _zz_when_ArraySlice_l118_25_1[5:0];
  assign _zz_when_ArraySlice_l173_25_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_25_1 = {1'd0, _zz_when_ArraySlice_l173_25_2};
  assign _zz_when_ArraySlice_l173_25_3 = (_zz_when_ArraySlice_l173_25_4 + _zz_when_ArraySlice_l173_25_9);
  assign _zz_when_ArraySlice_l173_25_4 = (_zz_when_ArraySlice_l173_25 - _zz_when_ArraySlice_l173_25_5);
  assign _zz_when_ArraySlice_l173_25_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_25_7);
  assign _zz_when_ArraySlice_l173_25_5 = {1'd0, _zz_when_ArraySlice_l173_25_6};
  assign _zz_when_ArraySlice_l173_25_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_25_7 = {2'd0, _zz_when_ArraySlice_l173_25_8};
  assign _zz_when_ArraySlice_l173_25_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_26 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_26_1);
  assign _zz_when_ArraySlice_l165_26_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_26_1 = {1'd0, _zz_when_ArraySlice_l165_26_2};
  assign _zz_when_ArraySlice_l166_26 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_26_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_26_2);
  assign _zz_when_ArraySlice_l166_26_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_26_3);
  assign _zz_when_ArraySlice_l166_26_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_26_3 = {1'd0, _zz_when_ArraySlice_l166_26_4};
  assign _zz__zz_when_ArraySlice_l112_26 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_26 = (_zz_when_ArraySlice_l113_26_1 - _zz_when_ArraySlice_l113_26_4);
  assign _zz_when_ArraySlice_l113_26_1 = (_zz_when_ArraySlice_l113_26_2 + _zz_when_ArraySlice_l113_26_3);
  assign _zz_when_ArraySlice_l113_26_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_26_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_26_4 = {1'd0, _zz_when_ArraySlice_l112_26};
  assign _zz__zz_when_ArraySlice_l173_26 = (_zz__zz_when_ArraySlice_l173_26_1 + _zz__zz_when_ArraySlice_l173_26_2);
  assign _zz__zz_when_ArraySlice_l173_26_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_26_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_26_3 = {1'd0, _zz_when_ArraySlice_l112_26};
  assign _zz_when_ArraySlice_l118_26_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_26 = _zz_when_ArraySlice_l118_26_1[5:0];
  assign _zz_when_ArraySlice_l173_26_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_26_1 = {1'd0, _zz_when_ArraySlice_l173_26_2};
  assign _zz_when_ArraySlice_l173_26_3 = (_zz_when_ArraySlice_l173_26_4 + _zz_when_ArraySlice_l173_26_9);
  assign _zz_when_ArraySlice_l173_26_4 = (_zz_when_ArraySlice_l173_26 - _zz_when_ArraySlice_l173_26_5);
  assign _zz_when_ArraySlice_l173_26_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_26_7);
  assign _zz_when_ArraySlice_l173_26_5 = {1'd0, _zz_when_ArraySlice_l173_26_6};
  assign _zz_when_ArraySlice_l173_26_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_26_7 = {1'd0, _zz_when_ArraySlice_l173_26_8};
  assign _zz_when_ArraySlice_l173_26_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_27 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_27_1);
  assign _zz_when_ArraySlice_l165_27_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_27_1 = {1'd0, _zz_when_ArraySlice_l165_27_2};
  assign _zz_when_ArraySlice_l166_27 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_27_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_27_2);
  assign _zz_when_ArraySlice_l166_27_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_27_3);
  assign _zz_when_ArraySlice_l166_27_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_27_3 = {1'd0, _zz_when_ArraySlice_l166_27_4};
  assign _zz__zz_when_ArraySlice_l112_27 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_27 = (_zz_when_ArraySlice_l113_27_1 - _zz_when_ArraySlice_l113_27_4);
  assign _zz_when_ArraySlice_l113_27_1 = (_zz_when_ArraySlice_l113_27_2 + _zz_when_ArraySlice_l113_27_3);
  assign _zz_when_ArraySlice_l113_27_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_27_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_27_4 = {1'd0, _zz_when_ArraySlice_l112_27};
  assign _zz__zz_when_ArraySlice_l173_27 = (_zz__zz_when_ArraySlice_l173_27_1 + _zz__zz_when_ArraySlice_l173_27_2);
  assign _zz__zz_when_ArraySlice_l173_27_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_27_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_27_3 = {1'd0, _zz_when_ArraySlice_l112_27};
  assign _zz_when_ArraySlice_l118_27_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_27 = _zz_when_ArraySlice_l118_27_1[5:0];
  assign _zz_when_ArraySlice_l173_27_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_27_1 = {1'd0, _zz_when_ArraySlice_l173_27_2};
  assign _zz_when_ArraySlice_l173_27_3 = (_zz_when_ArraySlice_l173_27_4 + _zz_when_ArraySlice_l173_27_9);
  assign _zz_when_ArraySlice_l173_27_4 = (_zz_when_ArraySlice_l173_27 - _zz_when_ArraySlice_l173_27_5);
  assign _zz_when_ArraySlice_l173_27_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_27_7);
  assign _zz_when_ArraySlice_l173_27_5 = {1'd0, _zz_when_ArraySlice_l173_27_6};
  assign _zz_when_ArraySlice_l173_27_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_27_7 = {1'd0, _zz_when_ArraySlice_l173_27_8};
  assign _zz_when_ArraySlice_l173_27_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_28 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_28_1);
  assign _zz_when_ArraySlice_l165_28_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_28 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_28_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_28_2);
  assign _zz_when_ArraySlice_l166_28_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_28_3);
  assign _zz_when_ArraySlice_l166_28_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_28 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_28 = (_zz_when_ArraySlice_l113_28_1 - _zz_when_ArraySlice_l113_28_4);
  assign _zz_when_ArraySlice_l113_28_1 = (_zz_when_ArraySlice_l113_28_2 + _zz_when_ArraySlice_l113_28_3);
  assign _zz_when_ArraySlice_l113_28_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_28_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_28_4 = {1'd0, _zz_when_ArraySlice_l112_28};
  assign _zz__zz_when_ArraySlice_l173_28 = (_zz__zz_when_ArraySlice_l173_28_1 + _zz__zz_when_ArraySlice_l173_28_2);
  assign _zz__zz_when_ArraySlice_l173_28_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_28_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_28_3 = {1'd0, _zz_when_ArraySlice_l112_28};
  assign _zz_when_ArraySlice_l118_28_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_28 = _zz_when_ArraySlice_l118_28_1[5:0];
  assign _zz_when_ArraySlice_l173_28_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_28_1 = {1'd0, _zz_when_ArraySlice_l173_28_2};
  assign _zz_when_ArraySlice_l173_28_3 = (_zz_when_ArraySlice_l173_28_4 + _zz_when_ArraySlice_l173_28_8);
  assign _zz_when_ArraySlice_l173_28_4 = (_zz_when_ArraySlice_l173_28 - _zz_when_ArraySlice_l173_28_5);
  assign _zz_when_ArraySlice_l173_28_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_28_7);
  assign _zz_when_ArraySlice_l173_28_5 = {1'd0, _zz_when_ArraySlice_l173_28_6};
  assign _zz_when_ArraySlice_l173_28_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_28_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_29 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_29_1);
  assign _zz_when_ArraySlice_l165_29_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_29_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_29 = {1'd0, _zz_when_ArraySlice_l166_29_1};
  assign _zz_when_ArraySlice_l166_29_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_29_3);
  assign _zz_when_ArraySlice_l166_29_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_29_4);
  assign _zz_when_ArraySlice_l166_29_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_29 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_29 = (_zz_when_ArraySlice_l113_29_1 - _zz_when_ArraySlice_l113_29_4);
  assign _zz_when_ArraySlice_l113_29_1 = (_zz_when_ArraySlice_l113_29_2 + _zz_when_ArraySlice_l113_29_3);
  assign _zz_when_ArraySlice_l113_29_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_29_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_29_4 = {1'd0, _zz_when_ArraySlice_l112_29};
  assign _zz__zz_when_ArraySlice_l173_29 = (_zz__zz_when_ArraySlice_l173_29_1 + _zz__zz_when_ArraySlice_l173_29_2);
  assign _zz__zz_when_ArraySlice_l173_29_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_29_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_29_3 = {1'd0, _zz_when_ArraySlice_l112_29};
  assign _zz_when_ArraySlice_l118_29_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_29 = _zz_when_ArraySlice_l118_29_1[5:0];
  assign _zz_when_ArraySlice_l173_29_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_29_1 = {2'd0, _zz_when_ArraySlice_l173_29_2};
  assign _zz_when_ArraySlice_l173_29_3 = (_zz_when_ArraySlice_l173_29_4 + _zz_when_ArraySlice_l173_29_8);
  assign _zz_when_ArraySlice_l173_29_4 = (_zz_when_ArraySlice_l173_29 - _zz_when_ArraySlice_l173_29_5);
  assign _zz_when_ArraySlice_l173_29_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_29_7);
  assign _zz_when_ArraySlice_l173_29_5 = {1'd0, _zz_when_ArraySlice_l173_29_6};
  assign _zz_when_ArraySlice_l173_29_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_29_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_30 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_30_1);
  assign _zz_when_ArraySlice_l165_30_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_30_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_30 = {1'd0, _zz_when_ArraySlice_l166_30_1};
  assign _zz_when_ArraySlice_l166_30_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_30_3);
  assign _zz_when_ArraySlice_l166_30_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_30_4);
  assign _zz_when_ArraySlice_l166_30_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_30 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_30 = (_zz_when_ArraySlice_l113_30_1 - _zz_when_ArraySlice_l113_30_4);
  assign _zz_when_ArraySlice_l113_30_1 = (_zz_when_ArraySlice_l113_30_2 + _zz_when_ArraySlice_l113_30_3);
  assign _zz_when_ArraySlice_l113_30_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_30_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_30_4 = {1'd0, _zz_when_ArraySlice_l112_30};
  assign _zz__zz_when_ArraySlice_l173_30 = (_zz__zz_when_ArraySlice_l173_30_1 + _zz__zz_when_ArraySlice_l173_30_2);
  assign _zz__zz_when_ArraySlice_l173_30_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_30_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_30_3 = {1'd0, _zz_when_ArraySlice_l112_30};
  assign _zz_when_ArraySlice_l118_30_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_30 = _zz_when_ArraySlice_l118_30_1[5:0];
  assign _zz_when_ArraySlice_l173_30_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_30_1 = {2'd0, _zz_when_ArraySlice_l173_30_2};
  assign _zz_when_ArraySlice_l173_30_3 = (_zz_when_ArraySlice_l173_30_4 + _zz_when_ArraySlice_l173_30_8);
  assign _zz_when_ArraySlice_l173_30_4 = (_zz_when_ArraySlice_l173_30 - _zz_when_ArraySlice_l173_30_5);
  assign _zz_when_ArraySlice_l173_30_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_30_7);
  assign _zz_when_ArraySlice_l173_30_5 = {1'd0, _zz_when_ArraySlice_l173_30_6};
  assign _zz_when_ArraySlice_l173_30_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_30_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_31 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_31_1);
  assign _zz_when_ArraySlice_l165_31_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_31_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_31 = {2'd0, _zz_when_ArraySlice_l166_31_1};
  assign _zz_when_ArraySlice_l166_31_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_31_3);
  assign _zz_when_ArraySlice_l166_31_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_31_4);
  assign _zz_when_ArraySlice_l166_31_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_31 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_31 = (_zz_when_ArraySlice_l113_31_1 - _zz_when_ArraySlice_l113_31_4);
  assign _zz_when_ArraySlice_l113_31_1 = (_zz_when_ArraySlice_l113_31_2 + _zz_when_ArraySlice_l113_31_3);
  assign _zz_when_ArraySlice_l113_31_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_31_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_31_4 = {1'd0, _zz_when_ArraySlice_l112_31};
  assign _zz__zz_when_ArraySlice_l173_31 = (_zz__zz_when_ArraySlice_l173_31_1 + _zz__zz_when_ArraySlice_l173_31_2);
  assign _zz__zz_when_ArraySlice_l173_31_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_31_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_31_3 = {1'd0, _zz_when_ArraySlice_l112_31};
  assign _zz_when_ArraySlice_l118_31_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_31 = _zz_when_ArraySlice_l118_31_1[5:0];
  assign _zz_when_ArraySlice_l173_31_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_31_1 = {3'd0, _zz_when_ArraySlice_l173_31_2};
  assign _zz_when_ArraySlice_l173_31_3 = (_zz_when_ArraySlice_l173_31_4 + _zz_when_ArraySlice_l173_31_8);
  assign _zz_when_ArraySlice_l173_31_4 = (_zz_when_ArraySlice_l173_31 - _zz_when_ArraySlice_l173_31_5);
  assign _zz_when_ArraySlice_l173_31_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_31_7);
  assign _zz_when_ArraySlice_l173_31_5 = {1'd0, _zz_when_ArraySlice_l173_31_6};
  assign _zz_when_ArraySlice_l173_31_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_31_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_0_31 = 1'b1;
  assign _zz_selectReadFifo_0_30 = {5'd0, _zz_selectReadFifo_0_31};
  assign _zz_when_ArraySlice_l448 = (_zz_when_ArraySlice_l448_1 % aReg);
  assign _zz_when_ArraySlice_l448_1 = (handshakeTimes_0_value + _zz_when_ArraySlice_l448_2);
  assign _zz_when_ArraySlice_l448_3 = 1'b1;
  assign _zz_when_ArraySlice_l448_2 = {12'd0, _zz_when_ArraySlice_l448_3};
  assign _zz_when_ArraySlice_l434 = (selectReadFifo_0 + _zz_when_ArraySlice_l434_1);
  assign _zz_when_ArraySlice_l434_2 = 3'b000;
  assign _zz_when_ArraySlice_l434_1 = {3'd0, _zz_when_ArraySlice_l434_2};
  assign _zz_when_ArraySlice_l455_1 = (_zz_when_ArraySlice_l455_2 - _zz_when_ArraySlice_l455_3);
  assign _zz_when_ArraySlice_l455 = {7'd0, _zz_when_ArraySlice_l455_1};
  assign _zz_when_ArraySlice_l455_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l455_4 = 1'b1;
  assign _zz_when_ArraySlice_l455_3 = {5'd0, _zz_when_ArraySlice_l455_4};
  assign _zz_when_ArraySlice_l373_1_1 = (selectReadFifo_1 + _zz_when_ArraySlice_l373_1_2);
  assign _zz_when_ArraySlice_l373_1_3 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l373_1_2 = {2'd0, _zz_when_ArraySlice_l373_1_3};
  assign _zz_when_ArraySlice_l374_1_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l374_1_3);
  assign _zz_when_ArraySlice_l374_1_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l374_1_3 = {2'd0, _zz_when_ArraySlice_l374_1_4};
  assign _zz__zz_outputStreamArrayData_1_valid_1 = (bReg * 1'b1);
  assign _zz__zz_outputStreamArrayData_1_valid = {2'd0, _zz__zz_outputStreamArrayData_1_valid_1};
  assign _zz_when_ArraySlice_l380_1_2 = 1'b1;
  assign _zz_when_ArraySlice_l380_1_1 = {6'd0, _zz_when_ArraySlice_l380_1_2};
  assign _zz_when_ArraySlice_l380_1_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l380_1_5);
  assign _zz_when_ArraySlice_l380_1_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l380_1_5 = {2'd0, _zz_when_ArraySlice_l380_1_6};
  assign _zz_when_ArraySlice_l381_1_2 = (_zz_when_ArraySlice_l381_1_3 - _zz_when_ArraySlice_l381_1_4);
  assign _zz_when_ArraySlice_l381_1_1 = {7'd0, _zz_when_ArraySlice_l381_1_2};
  assign _zz_when_ArraySlice_l381_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l381_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l381_1_4 = {5'd0, _zz_when_ArraySlice_l381_1_5};
  assign _zz_selectReadFifo_1 = (selectReadFifo_1 - _zz_selectReadFifo_1_1);
  assign _zz_selectReadFifo_1_1 = {3'd0, bReg};
  assign _zz_selectReadFifo_1_3 = 1'b1;
  assign _zz_selectReadFifo_1_2 = {5'd0, _zz_selectReadFifo_1_3};
  assign _zz_selectReadFifo_1_5 = 1'b1;
  assign _zz_selectReadFifo_1_4 = {5'd0, _zz_selectReadFifo_1_5};
  assign _zz_when_ArraySlice_l384_1_1 = (_zz_when_ArraySlice_l384_1_2 % aReg);
  assign _zz_when_ArraySlice_l384_1_2 = (handshakeTimes_1_value + _zz_when_ArraySlice_l384_1_3);
  assign _zz_when_ArraySlice_l384_1_4 = 1'b1;
  assign _zz_when_ArraySlice_l384_1_3 = {12'd0, _zz_when_ArraySlice_l384_1_4};
  assign _zz_when_ArraySlice_l389_1_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l389_1_3);
  assign _zz_when_ArraySlice_l389_1_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l389_1_3 = {2'd0, _zz_when_ArraySlice_l389_1_4};
  assign _zz_when_ArraySlice_l389_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l389_1_5 = {6'd0, _zz_when_ArraySlice_l389_1_6};
  assign _zz_when_ArraySlice_l390_1_2 = (_zz_when_ArraySlice_l390_1_3 - _zz_when_ArraySlice_l390_1_4);
  assign _zz_when_ArraySlice_l390_1_1 = {7'd0, _zz_when_ArraySlice_l390_1_2};
  assign _zz_when_ArraySlice_l390_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l390_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l390_1_4 = {5'd0, _zz_when_ArraySlice_l390_1_5};
  assign _zz__zz_when_ArraySlice_l94_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_3_1 = (_zz_when_ArraySlice_l95_3_2 - _zz_when_ArraySlice_l95_3_5);
  assign _zz_when_ArraySlice_l95_3_2 = (_zz_when_ArraySlice_l95_3_3 + _zz_when_ArraySlice_l95_3_4);
  assign _zz_when_ArraySlice_l95_3_3 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_3_4 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_3_5 = {1'd0, _zz_when_ArraySlice_l94_3};
  assign _zz__zz_when_ArraySlice_l392_1_1 = (_zz__zz_when_ArraySlice_l392_1_2 + _zz__zz_when_ArraySlice_l392_1_3);
  assign _zz__zz_when_ArraySlice_l392_1_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l392_1_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l392_1_4 = {1'd0, _zz_when_ArraySlice_l94_3};
  assign _zz_when_ArraySlice_l99_3_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_3 = _zz_when_ArraySlice_l99_3_1[5:0];
  assign _zz_when_ArraySlice_l392_1_1 = (outSliceNumb_1_value + _zz_when_ArraySlice_l392_1_2);
  assign _zz_when_ArraySlice_l392_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l392_1_2 = {6'd0, _zz_when_ArraySlice_l392_1_3};
  assign _zz_when_ArraySlice_l392_1_4 = (_zz_when_ArraySlice_l392_1 / aReg);
  assign _zz_selectReadFifo_1_6 = (selectReadFifo_1 - _zz_selectReadFifo_1_7);
  assign _zz_selectReadFifo_1_7 = {3'd0, bReg};
  assign _zz_selectReadFifo_1_9 = 1'b1;
  assign _zz_selectReadFifo_1_8 = {5'd0, _zz_selectReadFifo_1_9};
  assign _zz_selectReadFifo_1_10 = (selectReadFifo_1 + _zz_selectReadFifo_1_11);
  assign _zz_selectReadFifo_1_11 = (3'b111 * bReg);
  assign _zz_selectReadFifo_1_13 = 1'b1;
  assign _zz_selectReadFifo_1_12 = {5'd0, _zz_selectReadFifo_1_13};
  assign _zz_when_ArraySlice_l165_32 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_32_1);
  assign _zz_when_ArraySlice_l165_32_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_32_1 = {3'd0, _zz_when_ArraySlice_l165_32_2};
  assign _zz_when_ArraySlice_l166_32 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_32_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_32_3);
  assign _zz_when_ArraySlice_l166_32_1 = {1'd0, _zz_when_ArraySlice_l166_32_2};
  assign _zz_when_ArraySlice_l166_32_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_32_4);
  assign _zz_when_ArraySlice_l166_32_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_32_4 = {3'd0, _zz_when_ArraySlice_l166_32_5};
  assign _zz__zz_when_ArraySlice_l112_32 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_32 = (_zz_when_ArraySlice_l113_32_1 - _zz_when_ArraySlice_l113_32_4);
  assign _zz_when_ArraySlice_l113_32_1 = (_zz_when_ArraySlice_l113_32_2 + _zz_when_ArraySlice_l113_32_3);
  assign _zz_when_ArraySlice_l113_32_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_32_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_32_4 = {1'd0, _zz_when_ArraySlice_l112_32};
  assign _zz__zz_when_ArraySlice_l173_32 = (_zz__zz_when_ArraySlice_l173_32_1 + _zz__zz_when_ArraySlice_l173_32_2);
  assign _zz__zz_when_ArraySlice_l173_32_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_32_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_32_3 = {1'd0, _zz_when_ArraySlice_l112_32};
  assign _zz_when_ArraySlice_l118_32_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_32 = _zz_when_ArraySlice_l118_32_1[5:0];
  assign _zz_when_ArraySlice_l173_32_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_32_2 = (_zz_when_ArraySlice_l173_32_3 + _zz_when_ArraySlice_l173_32_8);
  assign _zz_when_ArraySlice_l173_32_3 = (_zz_when_ArraySlice_l173_32 - _zz_when_ArraySlice_l173_32_4);
  assign _zz_when_ArraySlice_l173_32_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_32_6);
  assign _zz_when_ArraySlice_l173_32_4 = {1'd0, _zz_when_ArraySlice_l173_32_5};
  assign _zz_when_ArraySlice_l173_32_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_32_6 = {3'd0, _zz_when_ArraySlice_l173_32_7};
  assign _zz_when_ArraySlice_l173_32_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_33 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_33_1);
  assign _zz_when_ArraySlice_l165_33_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_33_1 = {2'd0, _zz_when_ArraySlice_l165_33_2};
  assign _zz_when_ArraySlice_l166_33 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_33_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_33_2);
  assign _zz_when_ArraySlice_l166_33_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_33_3);
  assign _zz_when_ArraySlice_l166_33_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_33_3 = {2'd0, _zz_when_ArraySlice_l166_33_4};
  assign _zz__zz_when_ArraySlice_l112_33 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_33 = (_zz_when_ArraySlice_l113_33_1 - _zz_when_ArraySlice_l113_33_4);
  assign _zz_when_ArraySlice_l113_33_1 = (_zz_when_ArraySlice_l113_33_2 + _zz_when_ArraySlice_l113_33_3);
  assign _zz_when_ArraySlice_l113_33_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_33_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_33_4 = {1'd0, _zz_when_ArraySlice_l112_33};
  assign _zz__zz_when_ArraySlice_l173_33 = (_zz__zz_when_ArraySlice_l173_33_1 + _zz__zz_when_ArraySlice_l173_33_2);
  assign _zz__zz_when_ArraySlice_l173_33_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_33_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_33_3 = {1'd0, _zz_when_ArraySlice_l112_33};
  assign _zz_when_ArraySlice_l118_33_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_33 = _zz_when_ArraySlice_l118_33_1[5:0];
  assign _zz_when_ArraySlice_l173_33_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_33_1 = {1'd0, _zz_when_ArraySlice_l173_33_2};
  assign _zz_when_ArraySlice_l173_33_3 = (_zz_when_ArraySlice_l173_33_4 + _zz_when_ArraySlice_l173_33_9);
  assign _zz_when_ArraySlice_l173_33_4 = (_zz_when_ArraySlice_l173_33 - _zz_when_ArraySlice_l173_33_5);
  assign _zz_when_ArraySlice_l173_33_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_33_7);
  assign _zz_when_ArraySlice_l173_33_5 = {1'd0, _zz_when_ArraySlice_l173_33_6};
  assign _zz_when_ArraySlice_l173_33_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_33_7 = {2'd0, _zz_when_ArraySlice_l173_33_8};
  assign _zz_when_ArraySlice_l173_33_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_34 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_34_1);
  assign _zz_when_ArraySlice_l165_34_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_34_1 = {1'd0, _zz_when_ArraySlice_l165_34_2};
  assign _zz_when_ArraySlice_l166_34 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_34_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_34_2);
  assign _zz_when_ArraySlice_l166_34_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_34_3);
  assign _zz_when_ArraySlice_l166_34_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_34_3 = {1'd0, _zz_when_ArraySlice_l166_34_4};
  assign _zz__zz_when_ArraySlice_l112_34 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_34 = (_zz_when_ArraySlice_l113_34_1 - _zz_when_ArraySlice_l113_34_4);
  assign _zz_when_ArraySlice_l113_34_1 = (_zz_when_ArraySlice_l113_34_2 + _zz_when_ArraySlice_l113_34_3);
  assign _zz_when_ArraySlice_l113_34_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_34_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_34_4 = {1'd0, _zz_when_ArraySlice_l112_34};
  assign _zz__zz_when_ArraySlice_l173_34 = (_zz__zz_when_ArraySlice_l173_34_1 + _zz__zz_when_ArraySlice_l173_34_2);
  assign _zz__zz_when_ArraySlice_l173_34_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_34_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_34_3 = {1'd0, _zz_when_ArraySlice_l112_34};
  assign _zz_when_ArraySlice_l118_34_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_34 = _zz_when_ArraySlice_l118_34_1[5:0];
  assign _zz_when_ArraySlice_l173_34_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_34_1 = {1'd0, _zz_when_ArraySlice_l173_34_2};
  assign _zz_when_ArraySlice_l173_34_3 = (_zz_when_ArraySlice_l173_34_4 + _zz_when_ArraySlice_l173_34_9);
  assign _zz_when_ArraySlice_l173_34_4 = (_zz_when_ArraySlice_l173_34 - _zz_when_ArraySlice_l173_34_5);
  assign _zz_when_ArraySlice_l173_34_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_34_7);
  assign _zz_when_ArraySlice_l173_34_5 = {1'd0, _zz_when_ArraySlice_l173_34_6};
  assign _zz_when_ArraySlice_l173_34_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_34_7 = {1'd0, _zz_when_ArraySlice_l173_34_8};
  assign _zz_when_ArraySlice_l173_34_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_35 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_35_1);
  assign _zz_when_ArraySlice_l165_35_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_35_1 = {1'd0, _zz_when_ArraySlice_l165_35_2};
  assign _zz_when_ArraySlice_l166_35 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_35_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_35_2);
  assign _zz_when_ArraySlice_l166_35_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_35_3);
  assign _zz_when_ArraySlice_l166_35_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_35_3 = {1'd0, _zz_when_ArraySlice_l166_35_4};
  assign _zz__zz_when_ArraySlice_l112_35 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_35 = (_zz_when_ArraySlice_l113_35_1 - _zz_when_ArraySlice_l113_35_4);
  assign _zz_when_ArraySlice_l113_35_1 = (_zz_when_ArraySlice_l113_35_2 + _zz_when_ArraySlice_l113_35_3);
  assign _zz_when_ArraySlice_l113_35_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_35_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_35_4 = {1'd0, _zz_when_ArraySlice_l112_35};
  assign _zz__zz_when_ArraySlice_l173_35 = (_zz__zz_when_ArraySlice_l173_35_1 + _zz__zz_when_ArraySlice_l173_35_2);
  assign _zz__zz_when_ArraySlice_l173_35_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_35_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_35_3 = {1'd0, _zz_when_ArraySlice_l112_35};
  assign _zz_when_ArraySlice_l118_35_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_35 = _zz_when_ArraySlice_l118_35_1[5:0];
  assign _zz_when_ArraySlice_l173_35_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_35_1 = {1'd0, _zz_when_ArraySlice_l173_35_2};
  assign _zz_when_ArraySlice_l173_35_3 = (_zz_when_ArraySlice_l173_35_4 + _zz_when_ArraySlice_l173_35_9);
  assign _zz_when_ArraySlice_l173_35_4 = (_zz_when_ArraySlice_l173_35 - _zz_when_ArraySlice_l173_35_5);
  assign _zz_when_ArraySlice_l173_35_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_35_7);
  assign _zz_when_ArraySlice_l173_35_5 = {1'd0, _zz_when_ArraySlice_l173_35_6};
  assign _zz_when_ArraySlice_l173_35_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_35_7 = {1'd0, _zz_when_ArraySlice_l173_35_8};
  assign _zz_when_ArraySlice_l173_35_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_36 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_36_1);
  assign _zz_when_ArraySlice_l165_36_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_36 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_36_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_36_2);
  assign _zz_when_ArraySlice_l166_36_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_36_3);
  assign _zz_when_ArraySlice_l166_36_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_36 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_36 = (_zz_when_ArraySlice_l113_36_1 - _zz_when_ArraySlice_l113_36_4);
  assign _zz_when_ArraySlice_l113_36_1 = (_zz_when_ArraySlice_l113_36_2 + _zz_when_ArraySlice_l113_36_3);
  assign _zz_when_ArraySlice_l113_36_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_36_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_36_4 = {1'd0, _zz_when_ArraySlice_l112_36};
  assign _zz__zz_when_ArraySlice_l173_36 = (_zz__zz_when_ArraySlice_l173_36_1 + _zz__zz_when_ArraySlice_l173_36_2);
  assign _zz__zz_when_ArraySlice_l173_36_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_36_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_36_3 = {1'd0, _zz_when_ArraySlice_l112_36};
  assign _zz_when_ArraySlice_l118_36_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_36 = _zz_when_ArraySlice_l118_36_1[5:0];
  assign _zz_when_ArraySlice_l173_36_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_36_1 = {1'd0, _zz_when_ArraySlice_l173_36_2};
  assign _zz_when_ArraySlice_l173_36_3 = (_zz_when_ArraySlice_l173_36_4 + _zz_when_ArraySlice_l173_36_8);
  assign _zz_when_ArraySlice_l173_36_4 = (_zz_when_ArraySlice_l173_36 - _zz_when_ArraySlice_l173_36_5);
  assign _zz_when_ArraySlice_l173_36_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_36_7);
  assign _zz_when_ArraySlice_l173_36_5 = {1'd0, _zz_when_ArraySlice_l173_36_6};
  assign _zz_when_ArraySlice_l173_36_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_36_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_37 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_37_1);
  assign _zz_when_ArraySlice_l165_37_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_37_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_37 = {1'd0, _zz_when_ArraySlice_l166_37_1};
  assign _zz_when_ArraySlice_l166_37_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_37_3);
  assign _zz_when_ArraySlice_l166_37_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_37_4);
  assign _zz_when_ArraySlice_l166_37_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_37 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_37 = (_zz_when_ArraySlice_l113_37_1 - _zz_when_ArraySlice_l113_37_4);
  assign _zz_when_ArraySlice_l113_37_1 = (_zz_when_ArraySlice_l113_37_2 + _zz_when_ArraySlice_l113_37_3);
  assign _zz_when_ArraySlice_l113_37_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_37_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_37_4 = {1'd0, _zz_when_ArraySlice_l112_37};
  assign _zz__zz_when_ArraySlice_l173_37 = (_zz__zz_when_ArraySlice_l173_37_1 + _zz__zz_when_ArraySlice_l173_37_2);
  assign _zz__zz_when_ArraySlice_l173_37_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_37_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_37_3 = {1'd0, _zz_when_ArraySlice_l112_37};
  assign _zz_when_ArraySlice_l118_37_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_37 = _zz_when_ArraySlice_l118_37_1[5:0];
  assign _zz_when_ArraySlice_l173_37_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_37_1 = {2'd0, _zz_when_ArraySlice_l173_37_2};
  assign _zz_when_ArraySlice_l173_37_3 = (_zz_when_ArraySlice_l173_37_4 + _zz_when_ArraySlice_l173_37_8);
  assign _zz_when_ArraySlice_l173_37_4 = (_zz_when_ArraySlice_l173_37 - _zz_when_ArraySlice_l173_37_5);
  assign _zz_when_ArraySlice_l173_37_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_37_7);
  assign _zz_when_ArraySlice_l173_37_5 = {1'd0, _zz_when_ArraySlice_l173_37_6};
  assign _zz_when_ArraySlice_l173_37_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_37_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_38 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_38_1);
  assign _zz_when_ArraySlice_l165_38_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_38_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_38 = {1'd0, _zz_when_ArraySlice_l166_38_1};
  assign _zz_when_ArraySlice_l166_38_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_38_3);
  assign _zz_when_ArraySlice_l166_38_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_38_4);
  assign _zz_when_ArraySlice_l166_38_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_38 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_38 = (_zz_when_ArraySlice_l113_38_1 - _zz_when_ArraySlice_l113_38_4);
  assign _zz_when_ArraySlice_l113_38_1 = (_zz_when_ArraySlice_l113_38_2 + _zz_when_ArraySlice_l113_38_3);
  assign _zz_when_ArraySlice_l113_38_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_38_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_38_4 = {1'd0, _zz_when_ArraySlice_l112_38};
  assign _zz__zz_when_ArraySlice_l173_38 = (_zz__zz_when_ArraySlice_l173_38_1 + _zz__zz_when_ArraySlice_l173_38_2);
  assign _zz__zz_when_ArraySlice_l173_38_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_38_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_38_3 = {1'd0, _zz_when_ArraySlice_l112_38};
  assign _zz_when_ArraySlice_l118_38_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_38 = _zz_when_ArraySlice_l118_38_1[5:0];
  assign _zz_when_ArraySlice_l173_38_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_38_1 = {2'd0, _zz_when_ArraySlice_l173_38_2};
  assign _zz_when_ArraySlice_l173_38_3 = (_zz_when_ArraySlice_l173_38_4 + _zz_when_ArraySlice_l173_38_8);
  assign _zz_when_ArraySlice_l173_38_4 = (_zz_when_ArraySlice_l173_38 - _zz_when_ArraySlice_l173_38_5);
  assign _zz_when_ArraySlice_l173_38_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_38_7);
  assign _zz_when_ArraySlice_l173_38_5 = {1'd0, _zz_when_ArraySlice_l173_38_6};
  assign _zz_when_ArraySlice_l173_38_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_38_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_39 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_39_1);
  assign _zz_when_ArraySlice_l165_39_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_39_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_39 = {2'd0, _zz_when_ArraySlice_l166_39_1};
  assign _zz_when_ArraySlice_l166_39_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_39_3);
  assign _zz_when_ArraySlice_l166_39_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_39_4);
  assign _zz_when_ArraySlice_l166_39_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_39 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_39 = (_zz_when_ArraySlice_l113_39_1 - _zz_when_ArraySlice_l113_39_4);
  assign _zz_when_ArraySlice_l113_39_1 = (_zz_when_ArraySlice_l113_39_2 + _zz_when_ArraySlice_l113_39_3);
  assign _zz_when_ArraySlice_l113_39_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_39_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_39_4 = {1'd0, _zz_when_ArraySlice_l112_39};
  assign _zz__zz_when_ArraySlice_l173_39 = (_zz__zz_when_ArraySlice_l173_39_1 + _zz__zz_when_ArraySlice_l173_39_2);
  assign _zz__zz_when_ArraySlice_l173_39_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_39_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_39_3 = {1'd0, _zz_when_ArraySlice_l112_39};
  assign _zz_when_ArraySlice_l118_39_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_39 = _zz_when_ArraySlice_l118_39_1[5:0];
  assign _zz_when_ArraySlice_l173_39_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_39_1 = {3'd0, _zz_when_ArraySlice_l173_39_2};
  assign _zz_when_ArraySlice_l173_39_3 = (_zz_when_ArraySlice_l173_39_4 + _zz_when_ArraySlice_l173_39_8);
  assign _zz_when_ArraySlice_l173_39_4 = (_zz_when_ArraySlice_l173_39 - _zz_when_ArraySlice_l173_39_5);
  assign _zz_when_ArraySlice_l173_39_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_39_7);
  assign _zz_when_ArraySlice_l173_39_5 = {1'd0, _zz_when_ArraySlice_l173_39_6};
  assign _zz_when_ArraySlice_l173_39_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_39_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l401_1_1 = (_zz_when_ArraySlice_l401_1_2 + _zz_when_ArraySlice_l401_1_7);
  assign _zz_when_ArraySlice_l401_1_2 = (_zz_when_ArraySlice_l401_1_3 + _zz_when_ArraySlice_l401_1_5);
  assign _zz_when_ArraySlice_l401_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l401_1_4);
  assign _zz_when_ArraySlice_l401_1_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l401_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l401_1_5 = {5'd0, _zz_when_ArraySlice_l401_1_6};
  assign _zz_when_ArraySlice_l401_1_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l401_1_7 = {2'd0, _zz_when_ArraySlice_l401_1_8};
  assign _zz_selectReadFifo_1_15 = 1'b1;
  assign _zz_selectReadFifo_1_14 = {5'd0, _zz_selectReadFifo_1_15};
  assign _zz_when_ArraySlice_l405_1_1 = (_zz_when_ArraySlice_l405_1_2 % aReg);
  assign _zz_when_ArraySlice_l405_1_2 = (handshakeTimes_1_value + _zz_when_ArraySlice_l405_1_3);
  assign _zz_when_ArraySlice_l405_1_4 = 1'b1;
  assign _zz_when_ArraySlice_l405_1_3 = {12'd0, _zz_when_ArraySlice_l405_1_4};
  assign _zz_when_ArraySlice_l409_1_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l409_1_3);
  assign _zz_when_ArraySlice_l409_1_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l409_1_3 = {2'd0, _zz_when_ArraySlice_l409_1_4};
  assign _zz_when_ArraySlice_l410_1_2 = (_zz_when_ArraySlice_l410_1_3 - _zz_when_ArraySlice_l410_1_4);
  assign _zz_when_ArraySlice_l410_1_1 = {7'd0, _zz_when_ArraySlice_l410_1_2};
  assign _zz_when_ArraySlice_l410_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l410_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l410_1_4 = {5'd0, _zz_when_ArraySlice_l410_1_5};
  assign _zz__zz_when_ArraySlice_l94_4 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_4_1 = (_zz_when_ArraySlice_l95_4_2 - _zz_when_ArraySlice_l95_4_5);
  assign _zz_when_ArraySlice_l95_4_2 = (_zz_when_ArraySlice_l95_4_3 + _zz_when_ArraySlice_l95_4_4);
  assign _zz_when_ArraySlice_l95_4_3 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_4_4 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_4_5 = {1'd0, _zz_when_ArraySlice_l94_4};
  assign _zz__zz_when_ArraySlice_l412_1_1 = (_zz__zz_when_ArraySlice_l412_1_2 + _zz__zz_when_ArraySlice_l412_1_3);
  assign _zz__zz_when_ArraySlice_l412_1_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l412_1_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l412_1_4 = {1'd0, _zz_when_ArraySlice_l94_4};
  assign _zz_when_ArraySlice_l99_4_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_4 = _zz_when_ArraySlice_l99_4_1[5:0];
  assign _zz_when_ArraySlice_l412_1_1 = (outSliceNumb_1_value + _zz_when_ArraySlice_l412_1_2);
  assign _zz_when_ArraySlice_l412_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l412_1_2 = {6'd0, _zz_when_ArraySlice_l412_1_3};
  assign _zz_when_ArraySlice_l412_1_4 = (_zz_when_ArraySlice_l412_1 / aReg);
  assign _zz_selectReadFifo_1_16 = (selectReadFifo_1 - _zz_selectReadFifo_1_17);
  assign _zz_selectReadFifo_1_17 = {3'd0, bReg};
  assign _zz_selectReadFifo_1_19 = 1'b1;
  assign _zz_selectReadFifo_1_18 = {5'd0, _zz_selectReadFifo_1_19};
  assign _zz_selectReadFifo_1_20 = (selectReadFifo_1 + _zz_selectReadFifo_1_21);
  assign _zz_selectReadFifo_1_21 = (3'b111 * bReg);
  assign _zz_selectReadFifo_1_23 = 1'b1;
  assign _zz_selectReadFifo_1_22 = {5'd0, _zz_selectReadFifo_1_23};
  assign _zz_when_ArraySlice_l165_40 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_40_1);
  assign _zz_when_ArraySlice_l165_40_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_40_1 = {3'd0, _zz_when_ArraySlice_l165_40_2};
  assign _zz_when_ArraySlice_l166_40 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_40_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_40_3);
  assign _zz_when_ArraySlice_l166_40_1 = {1'd0, _zz_when_ArraySlice_l166_40_2};
  assign _zz_when_ArraySlice_l166_40_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_40_4);
  assign _zz_when_ArraySlice_l166_40_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_40_4 = {3'd0, _zz_when_ArraySlice_l166_40_5};
  assign _zz__zz_when_ArraySlice_l112_40 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_40 = (_zz_when_ArraySlice_l113_40_1 - _zz_when_ArraySlice_l113_40_4);
  assign _zz_when_ArraySlice_l113_40_1 = (_zz_when_ArraySlice_l113_40_2 + _zz_when_ArraySlice_l113_40_3);
  assign _zz_when_ArraySlice_l113_40_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_40_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_40_4 = {1'd0, _zz_when_ArraySlice_l112_40};
  assign _zz__zz_when_ArraySlice_l173_40 = (_zz__zz_when_ArraySlice_l173_40_1 + _zz__zz_when_ArraySlice_l173_40_2);
  assign _zz__zz_when_ArraySlice_l173_40_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_40_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_40_3 = {1'd0, _zz_when_ArraySlice_l112_40};
  assign _zz_when_ArraySlice_l118_40_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_40 = _zz_when_ArraySlice_l118_40_1[5:0];
  assign _zz_when_ArraySlice_l173_40_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_40_2 = (_zz_when_ArraySlice_l173_40_3 + _zz_when_ArraySlice_l173_40_8);
  assign _zz_when_ArraySlice_l173_40_3 = (_zz_when_ArraySlice_l173_40 - _zz_when_ArraySlice_l173_40_4);
  assign _zz_when_ArraySlice_l173_40_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_40_6);
  assign _zz_when_ArraySlice_l173_40_4 = {1'd0, _zz_when_ArraySlice_l173_40_5};
  assign _zz_when_ArraySlice_l173_40_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_40_6 = {3'd0, _zz_when_ArraySlice_l173_40_7};
  assign _zz_when_ArraySlice_l173_40_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_41 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_41_1);
  assign _zz_when_ArraySlice_l165_41_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_41_1 = {2'd0, _zz_when_ArraySlice_l165_41_2};
  assign _zz_when_ArraySlice_l166_41 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_41_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_41_2);
  assign _zz_when_ArraySlice_l166_41_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_41_3);
  assign _zz_when_ArraySlice_l166_41_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_41_3 = {2'd0, _zz_when_ArraySlice_l166_41_4};
  assign _zz__zz_when_ArraySlice_l112_41 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_41 = (_zz_when_ArraySlice_l113_41_1 - _zz_when_ArraySlice_l113_41_4);
  assign _zz_when_ArraySlice_l113_41_1 = (_zz_when_ArraySlice_l113_41_2 + _zz_when_ArraySlice_l113_41_3);
  assign _zz_when_ArraySlice_l113_41_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_41_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_41_4 = {1'd0, _zz_when_ArraySlice_l112_41};
  assign _zz__zz_when_ArraySlice_l173_41 = (_zz__zz_when_ArraySlice_l173_41_1 + _zz__zz_when_ArraySlice_l173_41_2);
  assign _zz__zz_when_ArraySlice_l173_41_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_41_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_41_3 = {1'd0, _zz_when_ArraySlice_l112_41};
  assign _zz_when_ArraySlice_l118_41_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_41 = _zz_when_ArraySlice_l118_41_1[5:0];
  assign _zz_when_ArraySlice_l173_41_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_41_1 = {1'd0, _zz_when_ArraySlice_l173_41_2};
  assign _zz_when_ArraySlice_l173_41_3 = (_zz_when_ArraySlice_l173_41_4 + _zz_when_ArraySlice_l173_41_9);
  assign _zz_when_ArraySlice_l173_41_4 = (_zz_when_ArraySlice_l173_41 - _zz_when_ArraySlice_l173_41_5);
  assign _zz_when_ArraySlice_l173_41_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_41_7);
  assign _zz_when_ArraySlice_l173_41_5 = {1'd0, _zz_when_ArraySlice_l173_41_6};
  assign _zz_when_ArraySlice_l173_41_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_41_7 = {2'd0, _zz_when_ArraySlice_l173_41_8};
  assign _zz_when_ArraySlice_l173_41_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_42 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_42_1);
  assign _zz_when_ArraySlice_l165_42_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_42_1 = {1'd0, _zz_when_ArraySlice_l165_42_2};
  assign _zz_when_ArraySlice_l166_42 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_42_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_42_2);
  assign _zz_when_ArraySlice_l166_42_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_42_3);
  assign _zz_when_ArraySlice_l166_42_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_42_3 = {1'd0, _zz_when_ArraySlice_l166_42_4};
  assign _zz__zz_when_ArraySlice_l112_42 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_42 = (_zz_when_ArraySlice_l113_42_1 - _zz_when_ArraySlice_l113_42_4);
  assign _zz_when_ArraySlice_l113_42_1 = (_zz_when_ArraySlice_l113_42_2 + _zz_when_ArraySlice_l113_42_3);
  assign _zz_when_ArraySlice_l113_42_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_42_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_42_4 = {1'd0, _zz_when_ArraySlice_l112_42};
  assign _zz__zz_when_ArraySlice_l173_42 = (_zz__zz_when_ArraySlice_l173_42_1 + _zz__zz_when_ArraySlice_l173_42_2);
  assign _zz__zz_when_ArraySlice_l173_42_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_42_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_42_3 = {1'd0, _zz_when_ArraySlice_l112_42};
  assign _zz_when_ArraySlice_l118_42_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_42 = _zz_when_ArraySlice_l118_42_1[5:0];
  assign _zz_when_ArraySlice_l173_42_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_42_1 = {1'd0, _zz_when_ArraySlice_l173_42_2};
  assign _zz_when_ArraySlice_l173_42_3 = (_zz_when_ArraySlice_l173_42_4 + _zz_when_ArraySlice_l173_42_9);
  assign _zz_when_ArraySlice_l173_42_4 = (_zz_when_ArraySlice_l173_42 - _zz_when_ArraySlice_l173_42_5);
  assign _zz_when_ArraySlice_l173_42_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_42_7);
  assign _zz_when_ArraySlice_l173_42_5 = {1'd0, _zz_when_ArraySlice_l173_42_6};
  assign _zz_when_ArraySlice_l173_42_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_42_7 = {1'd0, _zz_when_ArraySlice_l173_42_8};
  assign _zz_when_ArraySlice_l173_42_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_43 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_43_1);
  assign _zz_when_ArraySlice_l165_43_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_43_1 = {1'd0, _zz_when_ArraySlice_l165_43_2};
  assign _zz_when_ArraySlice_l166_43 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_43_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_43_2);
  assign _zz_when_ArraySlice_l166_43_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_43_3);
  assign _zz_when_ArraySlice_l166_43_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_43_3 = {1'd0, _zz_when_ArraySlice_l166_43_4};
  assign _zz__zz_when_ArraySlice_l112_43 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_43 = (_zz_when_ArraySlice_l113_43_1 - _zz_when_ArraySlice_l113_43_4);
  assign _zz_when_ArraySlice_l113_43_1 = (_zz_when_ArraySlice_l113_43_2 + _zz_when_ArraySlice_l113_43_3);
  assign _zz_when_ArraySlice_l113_43_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_43_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_43_4 = {1'd0, _zz_when_ArraySlice_l112_43};
  assign _zz__zz_when_ArraySlice_l173_43 = (_zz__zz_when_ArraySlice_l173_43_1 + _zz__zz_when_ArraySlice_l173_43_2);
  assign _zz__zz_when_ArraySlice_l173_43_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_43_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_43_3 = {1'd0, _zz_when_ArraySlice_l112_43};
  assign _zz_when_ArraySlice_l118_43_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_43 = _zz_when_ArraySlice_l118_43_1[5:0];
  assign _zz_when_ArraySlice_l173_43_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_43_1 = {1'd0, _zz_when_ArraySlice_l173_43_2};
  assign _zz_when_ArraySlice_l173_43_3 = (_zz_when_ArraySlice_l173_43_4 + _zz_when_ArraySlice_l173_43_9);
  assign _zz_when_ArraySlice_l173_43_4 = (_zz_when_ArraySlice_l173_43 - _zz_when_ArraySlice_l173_43_5);
  assign _zz_when_ArraySlice_l173_43_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_43_7);
  assign _zz_when_ArraySlice_l173_43_5 = {1'd0, _zz_when_ArraySlice_l173_43_6};
  assign _zz_when_ArraySlice_l173_43_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_43_7 = {1'd0, _zz_when_ArraySlice_l173_43_8};
  assign _zz_when_ArraySlice_l173_43_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_44 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_44_1);
  assign _zz_when_ArraySlice_l165_44_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_44 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_44_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_44_2);
  assign _zz_when_ArraySlice_l166_44_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_44_3);
  assign _zz_when_ArraySlice_l166_44_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_44 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_44 = (_zz_when_ArraySlice_l113_44_1 - _zz_when_ArraySlice_l113_44_4);
  assign _zz_when_ArraySlice_l113_44_1 = (_zz_when_ArraySlice_l113_44_2 + _zz_when_ArraySlice_l113_44_3);
  assign _zz_when_ArraySlice_l113_44_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_44_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_44_4 = {1'd0, _zz_when_ArraySlice_l112_44};
  assign _zz__zz_when_ArraySlice_l173_44 = (_zz__zz_when_ArraySlice_l173_44_1 + _zz__zz_when_ArraySlice_l173_44_2);
  assign _zz__zz_when_ArraySlice_l173_44_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_44_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_44_3 = {1'd0, _zz_when_ArraySlice_l112_44};
  assign _zz_when_ArraySlice_l118_44_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_44 = _zz_when_ArraySlice_l118_44_1[5:0];
  assign _zz_when_ArraySlice_l173_44_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_44_1 = {1'd0, _zz_when_ArraySlice_l173_44_2};
  assign _zz_when_ArraySlice_l173_44_3 = (_zz_when_ArraySlice_l173_44_4 + _zz_when_ArraySlice_l173_44_8);
  assign _zz_when_ArraySlice_l173_44_4 = (_zz_when_ArraySlice_l173_44 - _zz_when_ArraySlice_l173_44_5);
  assign _zz_when_ArraySlice_l173_44_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_44_7);
  assign _zz_when_ArraySlice_l173_44_5 = {1'd0, _zz_when_ArraySlice_l173_44_6};
  assign _zz_when_ArraySlice_l173_44_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_44_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_45 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_45_1);
  assign _zz_when_ArraySlice_l165_45_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_45_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_45 = {1'd0, _zz_when_ArraySlice_l166_45_1};
  assign _zz_when_ArraySlice_l166_45_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_45_3);
  assign _zz_when_ArraySlice_l166_45_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_45_4);
  assign _zz_when_ArraySlice_l166_45_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_45 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_45 = (_zz_when_ArraySlice_l113_45_1 - _zz_when_ArraySlice_l113_45_4);
  assign _zz_when_ArraySlice_l113_45_1 = (_zz_when_ArraySlice_l113_45_2 + _zz_when_ArraySlice_l113_45_3);
  assign _zz_when_ArraySlice_l113_45_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_45_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_45_4 = {1'd0, _zz_when_ArraySlice_l112_45};
  assign _zz__zz_when_ArraySlice_l173_45 = (_zz__zz_when_ArraySlice_l173_45_1 + _zz__zz_when_ArraySlice_l173_45_2);
  assign _zz__zz_when_ArraySlice_l173_45_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_45_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_45_3 = {1'd0, _zz_when_ArraySlice_l112_45};
  assign _zz_when_ArraySlice_l118_45_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_45 = _zz_when_ArraySlice_l118_45_1[5:0];
  assign _zz_when_ArraySlice_l173_45_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_45_1 = {2'd0, _zz_when_ArraySlice_l173_45_2};
  assign _zz_when_ArraySlice_l173_45_3 = (_zz_when_ArraySlice_l173_45_4 + _zz_when_ArraySlice_l173_45_8);
  assign _zz_when_ArraySlice_l173_45_4 = (_zz_when_ArraySlice_l173_45 - _zz_when_ArraySlice_l173_45_5);
  assign _zz_when_ArraySlice_l173_45_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_45_7);
  assign _zz_when_ArraySlice_l173_45_5 = {1'd0, _zz_when_ArraySlice_l173_45_6};
  assign _zz_when_ArraySlice_l173_45_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_45_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_46 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_46_1);
  assign _zz_when_ArraySlice_l165_46_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_46_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_46 = {1'd0, _zz_when_ArraySlice_l166_46_1};
  assign _zz_when_ArraySlice_l166_46_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_46_3);
  assign _zz_when_ArraySlice_l166_46_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_46_4);
  assign _zz_when_ArraySlice_l166_46_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_46 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_46 = (_zz_when_ArraySlice_l113_46_1 - _zz_when_ArraySlice_l113_46_4);
  assign _zz_when_ArraySlice_l113_46_1 = (_zz_when_ArraySlice_l113_46_2 + _zz_when_ArraySlice_l113_46_3);
  assign _zz_when_ArraySlice_l113_46_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_46_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_46_4 = {1'd0, _zz_when_ArraySlice_l112_46};
  assign _zz__zz_when_ArraySlice_l173_46 = (_zz__zz_when_ArraySlice_l173_46_1 + _zz__zz_when_ArraySlice_l173_46_2);
  assign _zz__zz_when_ArraySlice_l173_46_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_46_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_46_3 = {1'd0, _zz_when_ArraySlice_l112_46};
  assign _zz_when_ArraySlice_l118_46_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_46 = _zz_when_ArraySlice_l118_46_1[5:0];
  assign _zz_when_ArraySlice_l173_46_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_46_1 = {2'd0, _zz_when_ArraySlice_l173_46_2};
  assign _zz_when_ArraySlice_l173_46_3 = (_zz_when_ArraySlice_l173_46_4 + _zz_when_ArraySlice_l173_46_8);
  assign _zz_when_ArraySlice_l173_46_4 = (_zz_when_ArraySlice_l173_46 - _zz_when_ArraySlice_l173_46_5);
  assign _zz_when_ArraySlice_l173_46_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_46_7);
  assign _zz_when_ArraySlice_l173_46_5 = {1'd0, _zz_when_ArraySlice_l173_46_6};
  assign _zz_when_ArraySlice_l173_46_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_46_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_47 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_47_1);
  assign _zz_when_ArraySlice_l165_47_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_47_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_47 = {2'd0, _zz_when_ArraySlice_l166_47_1};
  assign _zz_when_ArraySlice_l166_47_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_47_3);
  assign _zz_when_ArraySlice_l166_47_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_47_4);
  assign _zz_when_ArraySlice_l166_47_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_47 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_47 = (_zz_when_ArraySlice_l113_47_1 - _zz_when_ArraySlice_l113_47_4);
  assign _zz_when_ArraySlice_l113_47_1 = (_zz_when_ArraySlice_l113_47_2 + _zz_when_ArraySlice_l113_47_3);
  assign _zz_when_ArraySlice_l113_47_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_47_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_47_4 = {1'd0, _zz_when_ArraySlice_l112_47};
  assign _zz__zz_when_ArraySlice_l173_47 = (_zz__zz_when_ArraySlice_l173_47_1 + _zz__zz_when_ArraySlice_l173_47_2);
  assign _zz__zz_when_ArraySlice_l173_47_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_47_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_47_3 = {1'd0, _zz_when_ArraySlice_l112_47};
  assign _zz_when_ArraySlice_l118_47_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_47 = _zz_when_ArraySlice_l118_47_1[5:0];
  assign _zz_when_ArraySlice_l173_47_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_47_1 = {3'd0, _zz_when_ArraySlice_l173_47_2};
  assign _zz_when_ArraySlice_l173_47_3 = (_zz_when_ArraySlice_l173_47_4 + _zz_when_ArraySlice_l173_47_8);
  assign _zz_when_ArraySlice_l173_47_4 = (_zz_when_ArraySlice_l173_47 - _zz_when_ArraySlice_l173_47_5);
  assign _zz_when_ArraySlice_l173_47_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_47_7);
  assign _zz_when_ArraySlice_l173_47_5 = {1'd0, _zz_when_ArraySlice_l173_47_6};
  assign _zz_when_ArraySlice_l173_47_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_47_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l421_1_1 = (_zz_when_ArraySlice_l421_1_2 + _zz_when_ArraySlice_l421_1_7);
  assign _zz_when_ArraySlice_l421_1_2 = (_zz_when_ArraySlice_l421_1_3 + _zz_when_ArraySlice_l421_1_5);
  assign _zz_when_ArraySlice_l421_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l421_1_4);
  assign _zz_when_ArraySlice_l421_1_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l421_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l421_1_5 = {5'd0, _zz_when_ArraySlice_l421_1_6};
  assign _zz_when_ArraySlice_l421_1_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l421_1_7 = {2'd0, _zz_when_ArraySlice_l421_1_8};
  assign _zz_selectReadFifo_1_25 = 1'b1;
  assign _zz_selectReadFifo_1_24 = {5'd0, _zz_selectReadFifo_1_25};
  assign _zz_when_ArraySlice_l425_1_1 = (_zz_when_ArraySlice_l425_1_2 % aReg);
  assign _zz_when_ArraySlice_l425_1_2 = (handshakeTimes_1_value + _zz_when_ArraySlice_l425_1_3);
  assign _zz_when_ArraySlice_l425_1_4 = 1'b1;
  assign _zz_when_ArraySlice_l425_1_3 = {12'd0, _zz_when_ArraySlice_l425_1_4};
  assign _zz_when_ArraySlice_l436_1_2 = (_zz_when_ArraySlice_l436_1_3 - _zz_when_ArraySlice_l436_1_4);
  assign _zz_when_ArraySlice_l436_1_1 = {7'd0, _zz_when_ArraySlice_l436_1_2};
  assign _zz_when_ArraySlice_l436_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l436_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l436_1_4 = {5'd0, _zz_when_ArraySlice_l436_1_5};
  assign _zz__zz_when_ArraySlice_l94_5 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_5 = (_zz_when_ArraySlice_l95_5_1 - _zz_when_ArraySlice_l95_5_4);
  assign _zz_when_ArraySlice_l95_5_1 = (_zz_when_ArraySlice_l95_5_2 + _zz_when_ArraySlice_l95_5_3);
  assign _zz_when_ArraySlice_l95_5_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_5_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_5_4 = {1'd0, _zz_when_ArraySlice_l94_5};
  assign _zz__zz_when_ArraySlice_l437_1_1 = (_zz__zz_when_ArraySlice_l437_1_2 + _zz__zz_when_ArraySlice_l437_1_3);
  assign _zz__zz_when_ArraySlice_l437_1_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l437_1_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l437_1_4 = {1'd0, _zz_when_ArraySlice_l94_5};
  assign _zz_when_ArraySlice_l99_5_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_5 = _zz_when_ArraySlice_l99_5_1[5:0];
  assign _zz_when_ArraySlice_l437_1_1 = (outSliceNumb_1_value + _zz_when_ArraySlice_l437_1_2);
  assign _zz_when_ArraySlice_l437_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l437_1_2 = {6'd0, _zz_when_ArraySlice_l437_1_3};
  assign _zz_when_ArraySlice_l437_1_4 = (_zz_when_ArraySlice_l437_1 / aReg);
  assign _zz_selectReadFifo_1_26 = (selectReadFifo_1 - _zz_selectReadFifo_1_27);
  assign _zz_selectReadFifo_1_27 = {3'd0, bReg};
  assign _zz_selectReadFifo_1_29 = 1'b1;
  assign _zz_selectReadFifo_1_28 = {5'd0, _zz_selectReadFifo_1_29};
  assign _zz_when_ArraySlice_l165_48 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_48_1);
  assign _zz_when_ArraySlice_l165_48_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_48_1 = {3'd0, _zz_when_ArraySlice_l165_48_2};
  assign _zz_when_ArraySlice_l166_48 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_48_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_48_3);
  assign _zz_when_ArraySlice_l166_48_1 = {1'd0, _zz_when_ArraySlice_l166_48_2};
  assign _zz_when_ArraySlice_l166_48_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_48_4);
  assign _zz_when_ArraySlice_l166_48_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_48_4 = {3'd0, _zz_when_ArraySlice_l166_48_5};
  assign _zz__zz_when_ArraySlice_l112_48 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_48 = (_zz_when_ArraySlice_l113_48_1 - _zz_when_ArraySlice_l113_48_4);
  assign _zz_when_ArraySlice_l113_48_1 = (_zz_when_ArraySlice_l113_48_2 + _zz_when_ArraySlice_l113_48_3);
  assign _zz_when_ArraySlice_l113_48_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_48_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_48_4 = {1'd0, _zz_when_ArraySlice_l112_48};
  assign _zz__zz_when_ArraySlice_l173_48 = (_zz__zz_when_ArraySlice_l173_48_1 + _zz__zz_when_ArraySlice_l173_48_2);
  assign _zz__zz_when_ArraySlice_l173_48_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_48_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_48_3 = {1'd0, _zz_when_ArraySlice_l112_48};
  assign _zz_when_ArraySlice_l118_48_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_48 = _zz_when_ArraySlice_l118_48_1[5:0];
  assign _zz_when_ArraySlice_l173_48_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_48_2 = (_zz_when_ArraySlice_l173_48_3 + _zz_when_ArraySlice_l173_48_8);
  assign _zz_when_ArraySlice_l173_48_3 = (_zz_when_ArraySlice_l173_48 - _zz_when_ArraySlice_l173_48_4);
  assign _zz_when_ArraySlice_l173_48_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_48_6);
  assign _zz_when_ArraySlice_l173_48_4 = {1'd0, _zz_when_ArraySlice_l173_48_5};
  assign _zz_when_ArraySlice_l173_48_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_48_6 = {3'd0, _zz_when_ArraySlice_l173_48_7};
  assign _zz_when_ArraySlice_l173_48_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_49 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_49_1);
  assign _zz_when_ArraySlice_l165_49_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_49_1 = {2'd0, _zz_when_ArraySlice_l165_49_2};
  assign _zz_when_ArraySlice_l166_49 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_49_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_49_2);
  assign _zz_when_ArraySlice_l166_49_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_49_3);
  assign _zz_when_ArraySlice_l166_49_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_49_3 = {2'd0, _zz_when_ArraySlice_l166_49_4};
  assign _zz__zz_when_ArraySlice_l112_49 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_49 = (_zz_when_ArraySlice_l113_49_1 - _zz_when_ArraySlice_l113_49_4);
  assign _zz_when_ArraySlice_l113_49_1 = (_zz_when_ArraySlice_l113_49_2 + _zz_when_ArraySlice_l113_49_3);
  assign _zz_when_ArraySlice_l113_49_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_49_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_49_4 = {1'd0, _zz_when_ArraySlice_l112_49};
  assign _zz__zz_when_ArraySlice_l173_49 = (_zz__zz_when_ArraySlice_l173_49_1 + _zz__zz_when_ArraySlice_l173_49_2);
  assign _zz__zz_when_ArraySlice_l173_49_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_49_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_49_3 = {1'd0, _zz_when_ArraySlice_l112_49};
  assign _zz_when_ArraySlice_l118_49_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_49 = _zz_when_ArraySlice_l118_49_1[5:0];
  assign _zz_when_ArraySlice_l173_49_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_49_1 = {1'd0, _zz_when_ArraySlice_l173_49_2};
  assign _zz_when_ArraySlice_l173_49_3 = (_zz_when_ArraySlice_l173_49_4 + _zz_when_ArraySlice_l173_49_9);
  assign _zz_when_ArraySlice_l173_49_4 = (_zz_when_ArraySlice_l173_49 - _zz_when_ArraySlice_l173_49_5);
  assign _zz_when_ArraySlice_l173_49_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_49_7);
  assign _zz_when_ArraySlice_l173_49_5 = {1'd0, _zz_when_ArraySlice_l173_49_6};
  assign _zz_when_ArraySlice_l173_49_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_49_7 = {2'd0, _zz_when_ArraySlice_l173_49_8};
  assign _zz_when_ArraySlice_l173_49_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_50 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_50_1);
  assign _zz_when_ArraySlice_l165_50_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_50_1 = {1'd0, _zz_when_ArraySlice_l165_50_2};
  assign _zz_when_ArraySlice_l166_50 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_50_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_50_2);
  assign _zz_when_ArraySlice_l166_50_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_50_3);
  assign _zz_when_ArraySlice_l166_50_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_50_3 = {1'd0, _zz_when_ArraySlice_l166_50_4};
  assign _zz__zz_when_ArraySlice_l112_50 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_50 = (_zz_when_ArraySlice_l113_50_1 - _zz_when_ArraySlice_l113_50_4);
  assign _zz_when_ArraySlice_l113_50_1 = (_zz_when_ArraySlice_l113_50_2 + _zz_when_ArraySlice_l113_50_3);
  assign _zz_when_ArraySlice_l113_50_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_50_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_50_4 = {1'd0, _zz_when_ArraySlice_l112_50};
  assign _zz__zz_when_ArraySlice_l173_50 = (_zz__zz_when_ArraySlice_l173_50_1 + _zz__zz_when_ArraySlice_l173_50_2);
  assign _zz__zz_when_ArraySlice_l173_50_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_50_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_50_3 = {1'd0, _zz_when_ArraySlice_l112_50};
  assign _zz_when_ArraySlice_l118_50_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_50 = _zz_when_ArraySlice_l118_50_1[5:0];
  assign _zz_when_ArraySlice_l173_50_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_50_1 = {1'd0, _zz_when_ArraySlice_l173_50_2};
  assign _zz_when_ArraySlice_l173_50_3 = (_zz_when_ArraySlice_l173_50_4 + _zz_when_ArraySlice_l173_50_9);
  assign _zz_when_ArraySlice_l173_50_4 = (_zz_when_ArraySlice_l173_50 - _zz_when_ArraySlice_l173_50_5);
  assign _zz_when_ArraySlice_l173_50_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_50_7);
  assign _zz_when_ArraySlice_l173_50_5 = {1'd0, _zz_when_ArraySlice_l173_50_6};
  assign _zz_when_ArraySlice_l173_50_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_50_7 = {1'd0, _zz_when_ArraySlice_l173_50_8};
  assign _zz_when_ArraySlice_l173_50_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_51 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_51_1);
  assign _zz_when_ArraySlice_l165_51_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_51_1 = {1'd0, _zz_when_ArraySlice_l165_51_2};
  assign _zz_when_ArraySlice_l166_51 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_51_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_51_2);
  assign _zz_when_ArraySlice_l166_51_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_51_3);
  assign _zz_when_ArraySlice_l166_51_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_51_3 = {1'd0, _zz_when_ArraySlice_l166_51_4};
  assign _zz__zz_when_ArraySlice_l112_51 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_51 = (_zz_when_ArraySlice_l113_51_1 - _zz_when_ArraySlice_l113_51_4);
  assign _zz_when_ArraySlice_l113_51_1 = (_zz_when_ArraySlice_l113_51_2 + _zz_when_ArraySlice_l113_51_3);
  assign _zz_when_ArraySlice_l113_51_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_51_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_51_4 = {1'd0, _zz_when_ArraySlice_l112_51};
  assign _zz__zz_when_ArraySlice_l173_51 = (_zz__zz_when_ArraySlice_l173_51_1 + _zz__zz_when_ArraySlice_l173_51_2);
  assign _zz__zz_when_ArraySlice_l173_51_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_51_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_51_3 = {1'd0, _zz_when_ArraySlice_l112_51};
  assign _zz_when_ArraySlice_l118_51_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_51 = _zz_when_ArraySlice_l118_51_1[5:0];
  assign _zz_when_ArraySlice_l173_51_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_51_1 = {1'd0, _zz_when_ArraySlice_l173_51_2};
  assign _zz_when_ArraySlice_l173_51_3 = (_zz_when_ArraySlice_l173_51_4 + _zz_when_ArraySlice_l173_51_9);
  assign _zz_when_ArraySlice_l173_51_4 = (_zz_when_ArraySlice_l173_51 - _zz_when_ArraySlice_l173_51_5);
  assign _zz_when_ArraySlice_l173_51_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_51_7);
  assign _zz_when_ArraySlice_l173_51_5 = {1'd0, _zz_when_ArraySlice_l173_51_6};
  assign _zz_when_ArraySlice_l173_51_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_51_7 = {1'd0, _zz_when_ArraySlice_l173_51_8};
  assign _zz_when_ArraySlice_l173_51_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_52 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_52_1);
  assign _zz_when_ArraySlice_l165_52_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_52 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_52_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_52_2);
  assign _zz_when_ArraySlice_l166_52_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_52_3);
  assign _zz_when_ArraySlice_l166_52_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_52 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_52 = (_zz_when_ArraySlice_l113_52_1 - _zz_when_ArraySlice_l113_52_4);
  assign _zz_when_ArraySlice_l113_52_1 = (_zz_when_ArraySlice_l113_52_2 + _zz_when_ArraySlice_l113_52_3);
  assign _zz_when_ArraySlice_l113_52_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_52_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_52_4 = {1'd0, _zz_when_ArraySlice_l112_52};
  assign _zz__zz_when_ArraySlice_l173_52 = (_zz__zz_when_ArraySlice_l173_52_1 + _zz__zz_when_ArraySlice_l173_52_2);
  assign _zz__zz_when_ArraySlice_l173_52_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_52_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_52_3 = {1'd0, _zz_when_ArraySlice_l112_52};
  assign _zz_when_ArraySlice_l118_52_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_52 = _zz_when_ArraySlice_l118_52_1[5:0];
  assign _zz_when_ArraySlice_l173_52_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_52_1 = {1'd0, _zz_when_ArraySlice_l173_52_2};
  assign _zz_when_ArraySlice_l173_52_3 = (_zz_when_ArraySlice_l173_52_4 + _zz_when_ArraySlice_l173_52_8);
  assign _zz_when_ArraySlice_l173_52_4 = (_zz_when_ArraySlice_l173_52 - _zz_when_ArraySlice_l173_52_5);
  assign _zz_when_ArraySlice_l173_52_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_52_7);
  assign _zz_when_ArraySlice_l173_52_5 = {1'd0, _zz_when_ArraySlice_l173_52_6};
  assign _zz_when_ArraySlice_l173_52_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_52_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_53 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_53_1);
  assign _zz_when_ArraySlice_l165_53_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_53_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_53 = {1'd0, _zz_when_ArraySlice_l166_53_1};
  assign _zz_when_ArraySlice_l166_53_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_53_3);
  assign _zz_when_ArraySlice_l166_53_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_53_4);
  assign _zz_when_ArraySlice_l166_53_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_53 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_53 = (_zz_when_ArraySlice_l113_53_1 - _zz_when_ArraySlice_l113_53_4);
  assign _zz_when_ArraySlice_l113_53_1 = (_zz_when_ArraySlice_l113_53_2 + _zz_when_ArraySlice_l113_53_3);
  assign _zz_when_ArraySlice_l113_53_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_53_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_53_4 = {1'd0, _zz_when_ArraySlice_l112_53};
  assign _zz__zz_when_ArraySlice_l173_53 = (_zz__zz_when_ArraySlice_l173_53_1 + _zz__zz_when_ArraySlice_l173_53_2);
  assign _zz__zz_when_ArraySlice_l173_53_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_53_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_53_3 = {1'd0, _zz_when_ArraySlice_l112_53};
  assign _zz_when_ArraySlice_l118_53_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_53 = _zz_when_ArraySlice_l118_53_1[5:0];
  assign _zz_when_ArraySlice_l173_53_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_53_1 = {2'd0, _zz_when_ArraySlice_l173_53_2};
  assign _zz_when_ArraySlice_l173_53_3 = (_zz_when_ArraySlice_l173_53_4 + _zz_when_ArraySlice_l173_53_8);
  assign _zz_when_ArraySlice_l173_53_4 = (_zz_when_ArraySlice_l173_53 - _zz_when_ArraySlice_l173_53_5);
  assign _zz_when_ArraySlice_l173_53_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_53_7);
  assign _zz_when_ArraySlice_l173_53_5 = {1'd0, _zz_when_ArraySlice_l173_53_6};
  assign _zz_when_ArraySlice_l173_53_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_53_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_54 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_54_1);
  assign _zz_when_ArraySlice_l165_54_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_54_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_54 = {1'd0, _zz_when_ArraySlice_l166_54_1};
  assign _zz_when_ArraySlice_l166_54_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_54_3);
  assign _zz_when_ArraySlice_l166_54_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_54_4);
  assign _zz_when_ArraySlice_l166_54_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_54 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_54 = (_zz_when_ArraySlice_l113_54_1 - _zz_when_ArraySlice_l113_54_4);
  assign _zz_when_ArraySlice_l113_54_1 = (_zz_when_ArraySlice_l113_54_2 + _zz_when_ArraySlice_l113_54_3);
  assign _zz_when_ArraySlice_l113_54_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_54_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_54_4 = {1'd0, _zz_when_ArraySlice_l112_54};
  assign _zz__zz_when_ArraySlice_l173_54 = (_zz__zz_when_ArraySlice_l173_54_1 + _zz__zz_when_ArraySlice_l173_54_2);
  assign _zz__zz_when_ArraySlice_l173_54_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_54_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_54_3 = {1'd0, _zz_when_ArraySlice_l112_54};
  assign _zz_when_ArraySlice_l118_54_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_54 = _zz_when_ArraySlice_l118_54_1[5:0];
  assign _zz_when_ArraySlice_l173_54_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_54_1 = {2'd0, _zz_when_ArraySlice_l173_54_2};
  assign _zz_when_ArraySlice_l173_54_3 = (_zz_when_ArraySlice_l173_54_4 + _zz_when_ArraySlice_l173_54_8);
  assign _zz_when_ArraySlice_l173_54_4 = (_zz_when_ArraySlice_l173_54 - _zz_when_ArraySlice_l173_54_5);
  assign _zz_when_ArraySlice_l173_54_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_54_7);
  assign _zz_when_ArraySlice_l173_54_5 = {1'd0, _zz_when_ArraySlice_l173_54_6};
  assign _zz_when_ArraySlice_l173_54_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_54_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_55 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_55_1);
  assign _zz_when_ArraySlice_l165_55_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_55_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_55 = {2'd0, _zz_when_ArraySlice_l166_55_1};
  assign _zz_when_ArraySlice_l166_55_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_55_3);
  assign _zz_when_ArraySlice_l166_55_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_55_4);
  assign _zz_when_ArraySlice_l166_55_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_55 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_55 = (_zz_when_ArraySlice_l113_55_1 - _zz_when_ArraySlice_l113_55_4);
  assign _zz_when_ArraySlice_l113_55_1 = (_zz_when_ArraySlice_l113_55_2 + _zz_when_ArraySlice_l113_55_3);
  assign _zz_when_ArraySlice_l113_55_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_55_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_55_4 = {1'd0, _zz_when_ArraySlice_l112_55};
  assign _zz__zz_when_ArraySlice_l173_55 = (_zz__zz_when_ArraySlice_l173_55_1 + _zz__zz_when_ArraySlice_l173_55_2);
  assign _zz__zz_when_ArraySlice_l173_55_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_55_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_55_3 = {1'd0, _zz_when_ArraySlice_l112_55};
  assign _zz_when_ArraySlice_l118_55_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_55 = _zz_when_ArraySlice_l118_55_1[5:0];
  assign _zz_when_ArraySlice_l173_55_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_55_1 = {3'd0, _zz_when_ArraySlice_l173_55_2};
  assign _zz_when_ArraySlice_l173_55_3 = (_zz_when_ArraySlice_l173_55_4 + _zz_when_ArraySlice_l173_55_8);
  assign _zz_when_ArraySlice_l173_55_4 = (_zz_when_ArraySlice_l173_55 - _zz_when_ArraySlice_l173_55_5);
  assign _zz_when_ArraySlice_l173_55_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_55_7);
  assign _zz_when_ArraySlice_l173_55_5 = {1'd0, _zz_when_ArraySlice_l173_55_6};
  assign _zz_when_ArraySlice_l173_55_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_55_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_1_31 = 1'b1;
  assign _zz_selectReadFifo_1_30 = {5'd0, _zz_selectReadFifo_1_31};
  assign _zz_when_ArraySlice_l448_1_1 = (_zz_when_ArraySlice_l448_1_2 % aReg);
  assign _zz_when_ArraySlice_l448_1_2 = (handshakeTimes_1_value + _zz_when_ArraySlice_l448_1_3);
  assign _zz_when_ArraySlice_l448_1_4 = 1'b1;
  assign _zz_when_ArraySlice_l448_1_3 = {12'd0, _zz_when_ArraySlice_l448_1_4};
  assign _zz_when_ArraySlice_l434_1_1 = (selectReadFifo_1 + _zz_when_ArraySlice_l434_1_2);
  assign _zz_when_ArraySlice_l434_1_3 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l434_1_2 = {2'd0, _zz_when_ArraySlice_l434_1_3};
  assign _zz_when_ArraySlice_l455_1_2 = (_zz_when_ArraySlice_l455_1_3 - _zz_when_ArraySlice_l455_1_4);
  assign _zz_when_ArraySlice_l455_1_1 = {7'd0, _zz_when_ArraySlice_l455_1_2};
  assign _zz_when_ArraySlice_l455_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l455_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l455_1_4 = {5'd0, _zz_when_ArraySlice_l455_1_5};
  assign _zz_when_ArraySlice_l373_2_1 = (selectReadFifo_2 + _zz_when_ArraySlice_l373_2_2);
  assign _zz_when_ArraySlice_l373_2_3 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l373_2_2 = {1'd0, _zz_when_ArraySlice_l373_2_3};
  assign _zz_when_ArraySlice_l374_2_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l374_2_3);
  assign _zz_when_ArraySlice_l374_2_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l374_2_3 = {1'd0, _zz_when_ArraySlice_l374_2_4};
  assign _zz__zz_outputStreamArrayData_2_valid_1 = (bReg * 2'b10);
  assign _zz__zz_outputStreamArrayData_2_valid = {1'd0, _zz__zz_outputStreamArrayData_2_valid_1};
  assign _zz_when_ArraySlice_l380_2_2 = 1'b1;
  assign _zz_when_ArraySlice_l380_2_1 = {6'd0, _zz_when_ArraySlice_l380_2_2};
  assign _zz_when_ArraySlice_l380_2_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l380_2_5);
  assign _zz_when_ArraySlice_l380_2_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l380_2_5 = {1'd0, _zz_when_ArraySlice_l380_2_6};
  assign _zz_when_ArraySlice_l381_2_2 = (_zz_when_ArraySlice_l381_2_3 - _zz_when_ArraySlice_l381_2_4);
  assign _zz_when_ArraySlice_l381_2_1 = {7'd0, _zz_when_ArraySlice_l381_2_2};
  assign _zz_when_ArraySlice_l381_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l381_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l381_2_4 = {5'd0, _zz_when_ArraySlice_l381_2_5};
  assign _zz_selectReadFifo_2 = (selectReadFifo_2 - _zz_selectReadFifo_2_1);
  assign _zz_selectReadFifo_2_1 = {3'd0, bReg};
  assign _zz_selectReadFifo_2_3 = 1'b1;
  assign _zz_selectReadFifo_2_2 = {5'd0, _zz_selectReadFifo_2_3};
  assign _zz_selectReadFifo_2_5 = 1'b1;
  assign _zz_selectReadFifo_2_4 = {5'd0, _zz_selectReadFifo_2_5};
  assign _zz_when_ArraySlice_l384_2_1 = (_zz_when_ArraySlice_l384_2_2 % aReg);
  assign _zz_when_ArraySlice_l384_2_2 = (handshakeTimes_2_value + _zz_when_ArraySlice_l384_2_3);
  assign _zz_when_ArraySlice_l384_2_4 = 1'b1;
  assign _zz_when_ArraySlice_l384_2_3 = {12'd0, _zz_when_ArraySlice_l384_2_4};
  assign _zz_when_ArraySlice_l389_2_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l389_2_3);
  assign _zz_when_ArraySlice_l389_2_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l389_2_3 = {1'd0, _zz_when_ArraySlice_l389_2_4};
  assign _zz_when_ArraySlice_l389_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l389_2_5 = {6'd0, _zz_when_ArraySlice_l389_2_6};
  assign _zz_when_ArraySlice_l390_2_2 = (_zz_when_ArraySlice_l390_2_3 - _zz_when_ArraySlice_l390_2_4);
  assign _zz_when_ArraySlice_l390_2_1 = {7'd0, _zz_when_ArraySlice_l390_2_2};
  assign _zz_when_ArraySlice_l390_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l390_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l390_2_4 = {5'd0, _zz_when_ArraySlice_l390_2_5};
  assign _zz__zz_when_ArraySlice_l94_6 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_6 = (_zz_when_ArraySlice_l95_6_1 - _zz_when_ArraySlice_l95_6_4);
  assign _zz_when_ArraySlice_l95_6_1 = (_zz_when_ArraySlice_l95_6_2 + _zz_when_ArraySlice_l95_6_3);
  assign _zz_when_ArraySlice_l95_6_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_6_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_6_4 = {1'd0, _zz_when_ArraySlice_l94_6};
  assign _zz__zz_when_ArraySlice_l392_2_1 = (_zz__zz_when_ArraySlice_l392_2_2 + _zz__zz_when_ArraySlice_l392_2_3);
  assign _zz__zz_when_ArraySlice_l392_2_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l392_2_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l392_2_4 = {1'd0, _zz_when_ArraySlice_l94_6};
  assign _zz_when_ArraySlice_l99_6_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_6 = _zz_when_ArraySlice_l99_6_1[5:0];
  assign _zz_when_ArraySlice_l392_2_1 = (outSliceNumb_2_value + _zz_when_ArraySlice_l392_2_2);
  assign _zz_when_ArraySlice_l392_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l392_2_2 = {6'd0, _zz_when_ArraySlice_l392_2_3};
  assign _zz_when_ArraySlice_l392_2_4 = (_zz_when_ArraySlice_l392_2 / aReg);
  assign _zz_selectReadFifo_2_6 = (selectReadFifo_2 - _zz_selectReadFifo_2_7);
  assign _zz_selectReadFifo_2_7 = {3'd0, bReg};
  assign _zz_selectReadFifo_2_9 = 1'b1;
  assign _zz_selectReadFifo_2_8 = {5'd0, _zz_selectReadFifo_2_9};
  assign _zz_selectReadFifo_2_10 = (selectReadFifo_2 + _zz_selectReadFifo_2_11);
  assign _zz_selectReadFifo_2_11 = (3'b111 * bReg);
  assign _zz_selectReadFifo_2_13 = 1'b1;
  assign _zz_selectReadFifo_2_12 = {5'd0, _zz_selectReadFifo_2_13};
  assign _zz_when_ArraySlice_l165_56 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_56_1);
  assign _zz_when_ArraySlice_l165_56_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_56_1 = {3'd0, _zz_when_ArraySlice_l165_56_2};
  assign _zz_when_ArraySlice_l166_56 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_56_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_56_3);
  assign _zz_when_ArraySlice_l166_56_1 = {1'd0, _zz_when_ArraySlice_l166_56_2};
  assign _zz_when_ArraySlice_l166_56_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_56_4);
  assign _zz_when_ArraySlice_l166_56_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_56_4 = {3'd0, _zz_when_ArraySlice_l166_56_5};
  assign _zz__zz_when_ArraySlice_l112_56 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_56 = (_zz_when_ArraySlice_l113_56_1 - _zz_when_ArraySlice_l113_56_4);
  assign _zz_when_ArraySlice_l113_56_1 = (_zz_when_ArraySlice_l113_56_2 + _zz_when_ArraySlice_l113_56_3);
  assign _zz_when_ArraySlice_l113_56_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_56_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_56_4 = {1'd0, _zz_when_ArraySlice_l112_56};
  assign _zz__zz_when_ArraySlice_l173_56 = (_zz__zz_when_ArraySlice_l173_56_1 + _zz__zz_when_ArraySlice_l173_56_2);
  assign _zz__zz_when_ArraySlice_l173_56_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_56_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_56_3 = {1'd0, _zz_when_ArraySlice_l112_56};
  assign _zz_when_ArraySlice_l118_56_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_56 = _zz_when_ArraySlice_l118_56_1[5:0];
  assign _zz_when_ArraySlice_l173_56_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_56_2 = (_zz_when_ArraySlice_l173_56_3 + _zz_when_ArraySlice_l173_56_8);
  assign _zz_when_ArraySlice_l173_56_3 = (_zz_when_ArraySlice_l173_56 - _zz_when_ArraySlice_l173_56_4);
  assign _zz_when_ArraySlice_l173_56_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_56_6);
  assign _zz_when_ArraySlice_l173_56_4 = {1'd0, _zz_when_ArraySlice_l173_56_5};
  assign _zz_when_ArraySlice_l173_56_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_56_6 = {3'd0, _zz_when_ArraySlice_l173_56_7};
  assign _zz_when_ArraySlice_l173_56_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_57 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_57_1);
  assign _zz_when_ArraySlice_l165_57_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_57_1 = {2'd0, _zz_when_ArraySlice_l165_57_2};
  assign _zz_when_ArraySlice_l166_57 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_57_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_57_2);
  assign _zz_when_ArraySlice_l166_57_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_57_3);
  assign _zz_when_ArraySlice_l166_57_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_57_3 = {2'd0, _zz_when_ArraySlice_l166_57_4};
  assign _zz__zz_when_ArraySlice_l112_57 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_57 = (_zz_when_ArraySlice_l113_57_1 - _zz_when_ArraySlice_l113_57_4);
  assign _zz_when_ArraySlice_l113_57_1 = (_zz_when_ArraySlice_l113_57_2 + _zz_when_ArraySlice_l113_57_3);
  assign _zz_when_ArraySlice_l113_57_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_57_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_57_4 = {1'd0, _zz_when_ArraySlice_l112_57};
  assign _zz__zz_when_ArraySlice_l173_57 = (_zz__zz_when_ArraySlice_l173_57_1 + _zz__zz_when_ArraySlice_l173_57_2);
  assign _zz__zz_when_ArraySlice_l173_57_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_57_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_57_3 = {1'd0, _zz_when_ArraySlice_l112_57};
  assign _zz_when_ArraySlice_l118_57_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_57 = _zz_when_ArraySlice_l118_57_1[5:0];
  assign _zz_when_ArraySlice_l173_57_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_57_1 = {1'd0, _zz_when_ArraySlice_l173_57_2};
  assign _zz_when_ArraySlice_l173_57_3 = (_zz_when_ArraySlice_l173_57_4 + _zz_when_ArraySlice_l173_57_9);
  assign _zz_when_ArraySlice_l173_57_4 = (_zz_when_ArraySlice_l173_57 - _zz_when_ArraySlice_l173_57_5);
  assign _zz_when_ArraySlice_l173_57_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_57_7);
  assign _zz_when_ArraySlice_l173_57_5 = {1'd0, _zz_when_ArraySlice_l173_57_6};
  assign _zz_when_ArraySlice_l173_57_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_57_7 = {2'd0, _zz_when_ArraySlice_l173_57_8};
  assign _zz_when_ArraySlice_l173_57_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_58 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_58_1);
  assign _zz_when_ArraySlice_l165_58_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_58_1 = {1'd0, _zz_when_ArraySlice_l165_58_2};
  assign _zz_when_ArraySlice_l166_58 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_58_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_58_2);
  assign _zz_when_ArraySlice_l166_58_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_58_3);
  assign _zz_when_ArraySlice_l166_58_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_58_3 = {1'd0, _zz_when_ArraySlice_l166_58_4};
  assign _zz__zz_when_ArraySlice_l112_58 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_58 = (_zz_when_ArraySlice_l113_58_1 - _zz_when_ArraySlice_l113_58_4);
  assign _zz_when_ArraySlice_l113_58_1 = (_zz_when_ArraySlice_l113_58_2 + _zz_when_ArraySlice_l113_58_3);
  assign _zz_when_ArraySlice_l113_58_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_58_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_58_4 = {1'd0, _zz_when_ArraySlice_l112_58};
  assign _zz__zz_when_ArraySlice_l173_58 = (_zz__zz_when_ArraySlice_l173_58_1 + _zz__zz_when_ArraySlice_l173_58_2);
  assign _zz__zz_when_ArraySlice_l173_58_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_58_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_58_3 = {1'd0, _zz_when_ArraySlice_l112_58};
  assign _zz_when_ArraySlice_l118_58_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_58 = _zz_when_ArraySlice_l118_58_1[5:0];
  assign _zz_when_ArraySlice_l173_58_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_58_1 = {1'd0, _zz_when_ArraySlice_l173_58_2};
  assign _zz_when_ArraySlice_l173_58_3 = (_zz_when_ArraySlice_l173_58_4 + _zz_when_ArraySlice_l173_58_9);
  assign _zz_when_ArraySlice_l173_58_4 = (_zz_when_ArraySlice_l173_58 - _zz_when_ArraySlice_l173_58_5);
  assign _zz_when_ArraySlice_l173_58_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_58_7);
  assign _zz_when_ArraySlice_l173_58_5 = {1'd0, _zz_when_ArraySlice_l173_58_6};
  assign _zz_when_ArraySlice_l173_58_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_58_7 = {1'd0, _zz_when_ArraySlice_l173_58_8};
  assign _zz_when_ArraySlice_l173_58_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_59 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_59_1);
  assign _zz_when_ArraySlice_l165_59_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_59_1 = {1'd0, _zz_when_ArraySlice_l165_59_2};
  assign _zz_when_ArraySlice_l166_59 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_59_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_59_2);
  assign _zz_when_ArraySlice_l166_59_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_59_3);
  assign _zz_when_ArraySlice_l166_59_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_59_3 = {1'd0, _zz_when_ArraySlice_l166_59_4};
  assign _zz__zz_when_ArraySlice_l112_59 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_59 = (_zz_when_ArraySlice_l113_59_1 - _zz_when_ArraySlice_l113_59_4);
  assign _zz_when_ArraySlice_l113_59_1 = (_zz_when_ArraySlice_l113_59_2 + _zz_when_ArraySlice_l113_59_3);
  assign _zz_when_ArraySlice_l113_59_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_59_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_59_4 = {1'd0, _zz_when_ArraySlice_l112_59};
  assign _zz__zz_when_ArraySlice_l173_59 = (_zz__zz_when_ArraySlice_l173_59_1 + _zz__zz_when_ArraySlice_l173_59_2);
  assign _zz__zz_when_ArraySlice_l173_59_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_59_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_59_3 = {1'd0, _zz_when_ArraySlice_l112_59};
  assign _zz_when_ArraySlice_l118_59_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_59 = _zz_when_ArraySlice_l118_59_1[5:0];
  assign _zz_when_ArraySlice_l173_59_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_59_1 = {1'd0, _zz_when_ArraySlice_l173_59_2};
  assign _zz_when_ArraySlice_l173_59_3 = (_zz_when_ArraySlice_l173_59_4 + _zz_when_ArraySlice_l173_59_9);
  assign _zz_when_ArraySlice_l173_59_4 = (_zz_when_ArraySlice_l173_59 - _zz_when_ArraySlice_l173_59_5);
  assign _zz_when_ArraySlice_l173_59_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_59_7);
  assign _zz_when_ArraySlice_l173_59_5 = {1'd0, _zz_when_ArraySlice_l173_59_6};
  assign _zz_when_ArraySlice_l173_59_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_59_7 = {1'd0, _zz_when_ArraySlice_l173_59_8};
  assign _zz_when_ArraySlice_l173_59_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_60 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_60_1);
  assign _zz_when_ArraySlice_l165_60_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_60 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_60_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_60_2);
  assign _zz_when_ArraySlice_l166_60_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_60_3);
  assign _zz_when_ArraySlice_l166_60_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_60 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_60 = (_zz_when_ArraySlice_l113_60_1 - _zz_when_ArraySlice_l113_60_4);
  assign _zz_when_ArraySlice_l113_60_1 = (_zz_when_ArraySlice_l113_60_2 + _zz_when_ArraySlice_l113_60_3);
  assign _zz_when_ArraySlice_l113_60_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_60_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_60_4 = {1'd0, _zz_when_ArraySlice_l112_60};
  assign _zz__zz_when_ArraySlice_l173_60 = (_zz__zz_when_ArraySlice_l173_60_1 + _zz__zz_when_ArraySlice_l173_60_2);
  assign _zz__zz_when_ArraySlice_l173_60_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_60_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_60_3 = {1'd0, _zz_when_ArraySlice_l112_60};
  assign _zz_when_ArraySlice_l118_60_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_60 = _zz_when_ArraySlice_l118_60_1[5:0];
  assign _zz_when_ArraySlice_l173_60_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_60_1 = {1'd0, _zz_when_ArraySlice_l173_60_2};
  assign _zz_when_ArraySlice_l173_60_3 = (_zz_when_ArraySlice_l173_60_4 + _zz_when_ArraySlice_l173_60_8);
  assign _zz_when_ArraySlice_l173_60_4 = (_zz_when_ArraySlice_l173_60 - _zz_when_ArraySlice_l173_60_5);
  assign _zz_when_ArraySlice_l173_60_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_60_7);
  assign _zz_when_ArraySlice_l173_60_5 = {1'd0, _zz_when_ArraySlice_l173_60_6};
  assign _zz_when_ArraySlice_l173_60_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_60_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_61 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_61_1);
  assign _zz_when_ArraySlice_l165_61_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_61_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_61 = {1'd0, _zz_when_ArraySlice_l166_61_1};
  assign _zz_when_ArraySlice_l166_61_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_61_3);
  assign _zz_when_ArraySlice_l166_61_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_61_4);
  assign _zz_when_ArraySlice_l166_61_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_61 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_61 = (_zz_when_ArraySlice_l113_61_1 - _zz_when_ArraySlice_l113_61_4);
  assign _zz_when_ArraySlice_l113_61_1 = (_zz_when_ArraySlice_l113_61_2 + _zz_when_ArraySlice_l113_61_3);
  assign _zz_when_ArraySlice_l113_61_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_61_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_61_4 = {1'd0, _zz_when_ArraySlice_l112_61};
  assign _zz__zz_when_ArraySlice_l173_61 = (_zz__zz_when_ArraySlice_l173_61_1 + _zz__zz_when_ArraySlice_l173_61_2);
  assign _zz__zz_when_ArraySlice_l173_61_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_61_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_61_3 = {1'd0, _zz_when_ArraySlice_l112_61};
  assign _zz_when_ArraySlice_l118_61_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_61 = _zz_when_ArraySlice_l118_61_1[5:0];
  assign _zz_when_ArraySlice_l173_61_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_61_1 = {2'd0, _zz_when_ArraySlice_l173_61_2};
  assign _zz_when_ArraySlice_l173_61_3 = (_zz_when_ArraySlice_l173_61_4 + _zz_when_ArraySlice_l173_61_8);
  assign _zz_when_ArraySlice_l173_61_4 = (_zz_when_ArraySlice_l173_61 - _zz_when_ArraySlice_l173_61_5);
  assign _zz_when_ArraySlice_l173_61_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_61_7);
  assign _zz_when_ArraySlice_l173_61_5 = {1'd0, _zz_when_ArraySlice_l173_61_6};
  assign _zz_when_ArraySlice_l173_61_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_61_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_62 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_62_1);
  assign _zz_when_ArraySlice_l165_62_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_62_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_62 = {1'd0, _zz_when_ArraySlice_l166_62_1};
  assign _zz_when_ArraySlice_l166_62_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_62_3);
  assign _zz_when_ArraySlice_l166_62_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_62_4);
  assign _zz_when_ArraySlice_l166_62_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_62 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_62 = (_zz_when_ArraySlice_l113_62_1 - _zz_when_ArraySlice_l113_62_4);
  assign _zz_when_ArraySlice_l113_62_1 = (_zz_when_ArraySlice_l113_62_2 + _zz_when_ArraySlice_l113_62_3);
  assign _zz_when_ArraySlice_l113_62_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_62_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_62_4 = {1'd0, _zz_when_ArraySlice_l112_62};
  assign _zz__zz_when_ArraySlice_l173_62 = (_zz__zz_when_ArraySlice_l173_62_1 + _zz__zz_when_ArraySlice_l173_62_2);
  assign _zz__zz_when_ArraySlice_l173_62_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_62_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_62_3 = {1'd0, _zz_when_ArraySlice_l112_62};
  assign _zz_when_ArraySlice_l118_62_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_62 = _zz_when_ArraySlice_l118_62_1[5:0];
  assign _zz_when_ArraySlice_l173_62_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_62_1 = {2'd0, _zz_when_ArraySlice_l173_62_2};
  assign _zz_when_ArraySlice_l173_62_3 = (_zz_when_ArraySlice_l173_62_4 + _zz_when_ArraySlice_l173_62_8);
  assign _zz_when_ArraySlice_l173_62_4 = (_zz_when_ArraySlice_l173_62 - _zz_when_ArraySlice_l173_62_5);
  assign _zz_when_ArraySlice_l173_62_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_62_7);
  assign _zz_when_ArraySlice_l173_62_5 = {1'd0, _zz_when_ArraySlice_l173_62_6};
  assign _zz_when_ArraySlice_l173_62_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_62_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_63 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_63_1);
  assign _zz_when_ArraySlice_l165_63_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_63_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_63 = {2'd0, _zz_when_ArraySlice_l166_63_1};
  assign _zz_when_ArraySlice_l166_63_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_63_3);
  assign _zz_when_ArraySlice_l166_63_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_63_4);
  assign _zz_when_ArraySlice_l166_63_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_63 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_63 = (_zz_when_ArraySlice_l113_63_1 - _zz_when_ArraySlice_l113_63_4);
  assign _zz_when_ArraySlice_l113_63_1 = (_zz_when_ArraySlice_l113_63_2 + _zz_when_ArraySlice_l113_63_3);
  assign _zz_when_ArraySlice_l113_63_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_63_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_63_4 = {1'd0, _zz_when_ArraySlice_l112_63};
  assign _zz__zz_when_ArraySlice_l173_63 = (_zz__zz_when_ArraySlice_l173_63_1 + _zz__zz_when_ArraySlice_l173_63_2);
  assign _zz__zz_when_ArraySlice_l173_63_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_63_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_63_3 = {1'd0, _zz_when_ArraySlice_l112_63};
  assign _zz_when_ArraySlice_l118_63_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_63 = _zz_when_ArraySlice_l118_63_1[5:0];
  assign _zz_when_ArraySlice_l173_63_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_63_1 = {3'd0, _zz_when_ArraySlice_l173_63_2};
  assign _zz_when_ArraySlice_l173_63_3 = (_zz_when_ArraySlice_l173_63_4 + _zz_when_ArraySlice_l173_63_8);
  assign _zz_when_ArraySlice_l173_63_4 = (_zz_when_ArraySlice_l173_63 - _zz_when_ArraySlice_l173_63_5);
  assign _zz_when_ArraySlice_l173_63_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_63_7);
  assign _zz_when_ArraySlice_l173_63_5 = {1'd0, _zz_when_ArraySlice_l173_63_6};
  assign _zz_when_ArraySlice_l173_63_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_63_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l401_2_1 = (_zz_when_ArraySlice_l401_2_2 + _zz_when_ArraySlice_l401_2_7);
  assign _zz_when_ArraySlice_l401_2_2 = (_zz_when_ArraySlice_l401_2_3 + _zz_when_ArraySlice_l401_2_5);
  assign _zz_when_ArraySlice_l401_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l401_2_4);
  assign _zz_when_ArraySlice_l401_2_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l401_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l401_2_5 = {5'd0, _zz_when_ArraySlice_l401_2_6};
  assign _zz_when_ArraySlice_l401_2_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l401_2_7 = {1'd0, _zz_when_ArraySlice_l401_2_8};
  assign _zz_selectReadFifo_2_15 = 1'b1;
  assign _zz_selectReadFifo_2_14 = {5'd0, _zz_selectReadFifo_2_15};
  assign _zz_when_ArraySlice_l405_2_1 = (_zz_when_ArraySlice_l405_2_2 % aReg);
  assign _zz_when_ArraySlice_l405_2_2 = (handshakeTimes_2_value + _zz_when_ArraySlice_l405_2_3);
  assign _zz_when_ArraySlice_l405_2_4 = 1'b1;
  assign _zz_when_ArraySlice_l405_2_3 = {12'd0, _zz_when_ArraySlice_l405_2_4};
  assign _zz_when_ArraySlice_l409_2_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l409_2_3);
  assign _zz_when_ArraySlice_l409_2_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l409_2_3 = {1'd0, _zz_when_ArraySlice_l409_2_4};
  assign _zz_when_ArraySlice_l410_2_2 = (_zz_when_ArraySlice_l410_2_3 - _zz_when_ArraySlice_l410_2_4);
  assign _zz_when_ArraySlice_l410_2_1 = {7'd0, _zz_when_ArraySlice_l410_2_2};
  assign _zz_when_ArraySlice_l410_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l410_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l410_2_4 = {5'd0, _zz_when_ArraySlice_l410_2_5};
  assign _zz__zz_when_ArraySlice_l94_7 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_7 = (_zz_when_ArraySlice_l95_7_1 - _zz_when_ArraySlice_l95_7_4);
  assign _zz_when_ArraySlice_l95_7_1 = (_zz_when_ArraySlice_l95_7_2 + _zz_when_ArraySlice_l95_7_3);
  assign _zz_when_ArraySlice_l95_7_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_7_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_7_4 = {1'd0, _zz_when_ArraySlice_l94_7};
  assign _zz__zz_when_ArraySlice_l412_2_1 = (_zz__zz_when_ArraySlice_l412_2_2 + _zz__zz_when_ArraySlice_l412_2_3);
  assign _zz__zz_when_ArraySlice_l412_2_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l412_2_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l412_2_4 = {1'd0, _zz_when_ArraySlice_l94_7};
  assign _zz_when_ArraySlice_l99_7_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_7 = _zz_when_ArraySlice_l99_7_1[5:0];
  assign _zz_when_ArraySlice_l412_2_1 = (outSliceNumb_2_value + _zz_when_ArraySlice_l412_2_2);
  assign _zz_when_ArraySlice_l412_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l412_2_2 = {6'd0, _zz_when_ArraySlice_l412_2_3};
  assign _zz_when_ArraySlice_l412_2_4 = (_zz_when_ArraySlice_l412_2 / aReg);
  assign _zz_selectReadFifo_2_16 = (selectReadFifo_2 - _zz_selectReadFifo_2_17);
  assign _zz_selectReadFifo_2_17 = {3'd0, bReg};
  assign _zz_selectReadFifo_2_19 = 1'b1;
  assign _zz_selectReadFifo_2_18 = {5'd0, _zz_selectReadFifo_2_19};
  assign _zz_selectReadFifo_2_20 = (selectReadFifo_2 + _zz_selectReadFifo_2_21);
  assign _zz_selectReadFifo_2_21 = (3'b111 * bReg);
  assign _zz_selectReadFifo_2_23 = 1'b1;
  assign _zz_selectReadFifo_2_22 = {5'd0, _zz_selectReadFifo_2_23};
  assign _zz_when_ArraySlice_l165_64 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_64_1);
  assign _zz_when_ArraySlice_l165_64_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_64_1 = {3'd0, _zz_when_ArraySlice_l165_64_2};
  assign _zz_when_ArraySlice_l166_64 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_64_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_64_3);
  assign _zz_when_ArraySlice_l166_64_1 = {1'd0, _zz_when_ArraySlice_l166_64_2};
  assign _zz_when_ArraySlice_l166_64_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_64_4);
  assign _zz_when_ArraySlice_l166_64_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_64_4 = {3'd0, _zz_when_ArraySlice_l166_64_5};
  assign _zz__zz_when_ArraySlice_l112_64 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_64 = (_zz_when_ArraySlice_l113_64_1 - _zz_when_ArraySlice_l113_64_4);
  assign _zz_when_ArraySlice_l113_64_1 = (_zz_when_ArraySlice_l113_64_2 + _zz_when_ArraySlice_l113_64_3);
  assign _zz_when_ArraySlice_l113_64_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_64_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_64_4 = {1'd0, _zz_when_ArraySlice_l112_64};
  assign _zz__zz_when_ArraySlice_l173_64 = (_zz__zz_when_ArraySlice_l173_64_1 + _zz__zz_when_ArraySlice_l173_64_2);
  assign _zz__zz_when_ArraySlice_l173_64_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_64_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_64_3 = {1'd0, _zz_when_ArraySlice_l112_64};
  assign _zz_when_ArraySlice_l118_64_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_64 = _zz_when_ArraySlice_l118_64_1[5:0];
  assign _zz_when_ArraySlice_l173_64_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_64_2 = (_zz_when_ArraySlice_l173_64_3 + _zz_when_ArraySlice_l173_64_8);
  assign _zz_when_ArraySlice_l173_64_3 = (_zz_when_ArraySlice_l173_64 - _zz_when_ArraySlice_l173_64_4);
  assign _zz_when_ArraySlice_l173_64_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_64_6);
  assign _zz_when_ArraySlice_l173_64_4 = {1'd0, _zz_when_ArraySlice_l173_64_5};
  assign _zz_when_ArraySlice_l173_64_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_64_6 = {3'd0, _zz_when_ArraySlice_l173_64_7};
  assign _zz_when_ArraySlice_l173_64_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_65 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_65_1);
  assign _zz_when_ArraySlice_l165_65_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_65_1 = {2'd0, _zz_when_ArraySlice_l165_65_2};
  assign _zz_when_ArraySlice_l166_65 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_65_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_65_2);
  assign _zz_when_ArraySlice_l166_65_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_65_3);
  assign _zz_when_ArraySlice_l166_65_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_65_3 = {2'd0, _zz_when_ArraySlice_l166_65_4};
  assign _zz__zz_when_ArraySlice_l112_65 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_65 = (_zz_when_ArraySlice_l113_65_1 - _zz_when_ArraySlice_l113_65_4);
  assign _zz_when_ArraySlice_l113_65_1 = (_zz_when_ArraySlice_l113_65_2 + _zz_when_ArraySlice_l113_65_3);
  assign _zz_when_ArraySlice_l113_65_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_65_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_65_4 = {1'd0, _zz_when_ArraySlice_l112_65};
  assign _zz__zz_when_ArraySlice_l173_65 = (_zz__zz_when_ArraySlice_l173_65_1 + _zz__zz_when_ArraySlice_l173_65_2);
  assign _zz__zz_when_ArraySlice_l173_65_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_65_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_65_3 = {1'd0, _zz_when_ArraySlice_l112_65};
  assign _zz_when_ArraySlice_l118_65_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_65 = _zz_when_ArraySlice_l118_65_1[5:0];
  assign _zz_when_ArraySlice_l173_65_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_65_1 = {1'd0, _zz_when_ArraySlice_l173_65_2};
  assign _zz_when_ArraySlice_l173_65_3 = (_zz_when_ArraySlice_l173_65_4 + _zz_when_ArraySlice_l173_65_9);
  assign _zz_when_ArraySlice_l173_65_4 = (_zz_when_ArraySlice_l173_65 - _zz_when_ArraySlice_l173_65_5);
  assign _zz_when_ArraySlice_l173_65_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_65_7);
  assign _zz_when_ArraySlice_l173_65_5 = {1'd0, _zz_when_ArraySlice_l173_65_6};
  assign _zz_when_ArraySlice_l173_65_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_65_7 = {2'd0, _zz_when_ArraySlice_l173_65_8};
  assign _zz_when_ArraySlice_l173_65_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_66 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_66_1);
  assign _zz_when_ArraySlice_l165_66_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_66_1 = {1'd0, _zz_when_ArraySlice_l165_66_2};
  assign _zz_when_ArraySlice_l166_66 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_66_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_66_2);
  assign _zz_when_ArraySlice_l166_66_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_66_3);
  assign _zz_when_ArraySlice_l166_66_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_66_3 = {1'd0, _zz_when_ArraySlice_l166_66_4};
  assign _zz__zz_when_ArraySlice_l112_66 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_66 = (_zz_when_ArraySlice_l113_66_1 - _zz_when_ArraySlice_l113_66_4);
  assign _zz_when_ArraySlice_l113_66_1 = (_zz_when_ArraySlice_l113_66_2 + _zz_when_ArraySlice_l113_66_3);
  assign _zz_when_ArraySlice_l113_66_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_66_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_66_4 = {1'd0, _zz_when_ArraySlice_l112_66};
  assign _zz__zz_when_ArraySlice_l173_66 = (_zz__zz_when_ArraySlice_l173_66_1 + _zz__zz_when_ArraySlice_l173_66_2);
  assign _zz__zz_when_ArraySlice_l173_66_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_66_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_66_3 = {1'd0, _zz_when_ArraySlice_l112_66};
  assign _zz_when_ArraySlice_l118_66_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_66 = _zz_when_ArraySlice_l118_66_1[5:0];
  assign _zz_when_ArraySlice_l173_66_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_66_1 = {1'd0, _zz_when_ArraySlice_l173_66_2};
  assign _zz_when_ArraySlice_l173_66_3 = (_zz_when_ArraySlice_l173_66_4 + _zz_when_ArraySlice_l173_66_9);
  assign _zz_when_ArraySlice_l173_66_4 = (_zz_when_ArraySlice_l173_66 - _zz_when_ArraySlice_l173_66_5);
  assign _zz_when_ArraySlice_l173_66_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_66_7);
  assign _zz_when_ArraySlice_l173_66_5 = {1'd0, _zz_when_ArraySlice_l173_66_6};
  assign _zz_when_ArraySlice_l173_66_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_66_7 = {1'd0, _zz_when_ArraySlice_l173_66_8};
  assign _zz_when_ArraySlice_l173_66_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_67 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_67_1);
  assign _zz_when_ArraySlice_l165_67_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_67_1 = {1'd0, _zz_when_ArraySlice_l165_67_2};
  assign _zz_when_ArraySlice_l166_67 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_67_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_67_2);
  assign _zz_when_ArraySlice_l166_67_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_67_3);
  assign _zz_when_ArraySlice_l166_67_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_67_3 = {1'd0, _zz_when_ArraySlice_l166_67_4};
  assign _zz__zz_when_ArraySlice_l112_67 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_67 = (_zz_when_ArraySlice_l113_67_1 - _zz_when_ArraySlice_l113_67_4);
  assign _zz_when_ArraySlice_l113_67_1 = (_zz_when_ArraySlice_l113_67_2 + _zz_when_ArraySlice_l113_67_3);
  assign _zz_when_ArraySlice_l113_67_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_67_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_67_4 = {1'd0, _zz_when_ArraySlice_l112_67};
  assign _zz__zz_when_ArraySlice_l173_67 = (_zz__zz_when_ArraySlice_l173_67_1 + _zz__zz_when_ArraySlice_l173_67_2);
  assign _zz__zz_when_ArraySlice_l173_67_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_67_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_67_3 = {1'd0, _zz_when_ArraySlice_l112_67};
  assign _zz_when_ArraySlice_l118_67_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_67 = _zz_when_ArraySlice_l118_67_1[5:0];
  assign _zz_when_ArraySlice_l173_67_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_67_1 = {1'd0, _zz_when_ArraySlice_l173_67_2};
  assign _zz_when_ArraySlice_l173_67_3 = (_zz_when_ArraySlice_l173_67_4 + _zz_when_ArraySlice_l173_67_9);
  assign _zz_when_ArraySlice_l173_67_4 = (_zz_when_ArraySlice_l173_67 - _zz_when_ArraySlice_l173_67_5);
  assign _zz_when_ArraySlice_l173_67_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_67_7);
  assign _zz_when_ArraySlice_l173_67_5 = {1'd0, _zz_when_ArraySlice_l173_67_6};
  assign _zz_when_ArraySlice_l173_67_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_67_7 = {1'd0, _zz_when_ArraySlice_l173_67_8};
  assign _zz_when_ArraySlice_l173_67_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_68 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_68_1);
  assign _zz_when_ArraySlice_l165_68_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_68 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_68_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_68_2);
  assign _zz_when_ArraySlice_l166_68_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_68_3);
  assign _zz_when_ArraySlice_l166_68_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_68 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_68 = (_zz_when_ArraySlice_l113_68_1 - _zz_when_ArraySlice_l113_68_4);
  assign _zz_when_ArraySlice_l113_68_1 = (_zz_when_ArraySlice_l113_68_2 + _zz_when_ArraySlice_l113_68_3);
  assign _zz_when_ArraySlice_l113_68_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_68_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_68_4 = {1'd0, _zz_when_ArraySlice_l112_68};
  assign _zz__zz_when_ArraySlice_l173_68 = (_zz__zz_when_ArraySlice_l173_68_1 + _zz__zz_when_ArraySlice_l173_68_2);
  assign _zz__zz_when_ArraySlice_l173_68_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_68_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_68_3 = {1'd0, _zz_when_ArraySlice_l112_68};
  assign _zz_when_ArraySlice_l118_68_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_68 = _zz_when_ArraySlice_l118_68_1[5:0];
  assign _zz_when_ArraySlice_l173_68_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_68_1 = {1'd0, _zz_when_ArraySlice_l173_68_2};
  assign _zz_when_ArraySlice_l173_68_3 = (_zz_when_ArraySlice_l173_68_4 + _zz_when_ArraySlice_l173_68_8);
  assign _zz_when_ArraySlice_l173_68_4 = (_zz_when_ArraySlice_l173_68 - _zz_when_ArraySlice_l173_68_5);
  assign _zz_when_ArraySlice_l173_68_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_68_7);
  assign _zz_when_ArraySlice_l173_68_5 = {1'd0, _zz_when_ArraySlice_l173_68_6};
  assign _zz_when_ArraySlice_l173_68_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_68_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_69 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_69_1);
  assign _zz_when_ArraySlice_l165_69_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_69_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_69 = {1'd0, _zz_when_ArraySlice_l166_69_1};
  assign _zz_when_ArraySlice_l166_69_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_69_3);
  assign _zz_when_ArraySlice_l166_69_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_69_4);
  assign _zz_when_ArraySlice_l166_69_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_69 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_69 = (_zz_when_ArraySlice_l113_69_1 - _zz_when_ArraySlice_l113_69_4);
  assign _zz_when_ArraySlice_l113_69_1 = (_zz_when_ArraySlice_l113_69_2 + _zz_when_ArraySlice_l113_69_3);
  assign _zz_when_ArraySlice_l113_69_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_69_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_69_4 = {1'd0, _zz_when_ArraySlice_l112_69};
  assign _zz__zz_when_ArraySlice_l173_69 = (_zz__zz_when_ArraySlice_l173_69_1 + _zz__zz_when_ArraySlice_l173_69_2);
  assign _zz__zz_when_ArraySlice_l173_69_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_69_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_69_3 = {1'd0, _zz_when_ArraySlice_l112_69};
  assign _zz_when_ArraySlice_l118_69_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_69 = _zz_when_ArraySlice_l118_69_1[5:0];
  assign _zz_when_ArraySlice_l173_69_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_69_1 = {2'd0, _zz_when_ArraySlice_l173_69_2};
  assign _zz_when_ArraySlice_l173_69_3 = (_zz_when_ArraySlice_l173_69_4 + _zz_when_ArraySlice_l173_69_8);
  assign _zz_when_ArraySlice_l173_69_4 = (_zz_when_ArraySlice_l173_69 - _zz_when_ArraySlice_l173_69_5);
  assign _zz_when_ArraySlice_l173_69_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_69_7);
  assign _zz_when_ArraySlice_l173_69_5 = {1'd0, _zz_when_ArraySlice_l173_69_6};
  assign _zz_when_ArraySlice_l173_69_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_69_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_70 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_70_1);
  assign _zz_when_ArraySlice_l165_70_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_70_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_70 = {1'd0, _zz_when_ArraySlice_l166_70_1};
  assign _zz_when_ArraySlice_l166_70_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_70_3);
  assign _zz_when_ArraySlice_l166_70_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_70_4);
  assign _zz_when_ArraySlice_l166_70_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_70 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_70 = (_zz_when_ArraySlice_l113_70_1 - _zz_when_ArraySlice_l113_70_4);
  assign _zz_when_ArraySlice_l113_70_1 = (_zz_when_ArraySlice_l113_70_2 + _zz_when_ArraySlice_l113_70_3);
  assign _zz_when_ArraySlice_l113_70_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_70_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_70_4 = {1'd0, _zz_when_ArraySlice_l112_70};
  assign _zz__zz_when_ArraySlice_l173_70 = (_zz__zz_when_ArraySlice_l173_70_1 + _zz__zz_when_ArraySlice_l173_70_2);
  assign _zz__zz_when_ArraySlice_l173_70_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_70_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_70_3 = {1'd0, _zz_when_ArraySlice_l112_70};
  assign _zz_when_ArraySlice_l118_70_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_70 = _zz_when_ArraySlice_l118_70_1[5:0];
  assign _zz_when_ArraySlice_l173_70_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_70_1 = {2'd0, _zz_when_ArraySlice_l173_70_2};
  assign _zz_when_ArraySlice_l173_70_3 = (_zz_when_ArraySlice_l173_70_4 + _zz_when_ArraySlice_l173_70_8);
  assign _zz_when_ArraySlice_l173_70_4 = (_zz_when_ArraySlice_l173_70 - _zz_when_ArraySlice_l173_70_5);
  assign _zz_when_ArraySlice_l173_70_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_70_7);
  assign _zz_when_ArraySlice_l173_70_5 = {1'd0, _zz_when_ArraySlice_l173_70_6};
  assign _zz_when_ArraySlice_l173_70_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_70_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_71 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_71_1);
  assign _zz_when_ArraySlice_l165_71_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_71_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_71 = {2'd0, _zz_when_ArraySlice_l166_71_1};
  assign _zz_when_ArraySlice_l166_71_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_71_3);
  assign _zz_when_ArraySlice_l166_71_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_71_4);
  assign _zz_when_ArraySlice_l166_71_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_71 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_71 = (_zz_when_ArraySlice_l113_71_1 - _zz_when_ArraySlice_l113_71_4);
  assign _zz_when_ArraySlice_l113_71_1 = (_zz_when_ArraySlice_l113_71_2 + _zz_when_ArraySlice_l113_71_3);
  assign _zz_when_ArraySlice_l113_71_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_71_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_71_4 = {1'd0, _zz_when_ArraySlice_l112_71};
  assign _zz__zz_when_ArraySlice_l173_71 = (_zz__zz_when_ArraySlice_l173_71_1 + _zz__zz_when_ArraySlice_l173_71_2);
  assign _zz__zz_when_ArraySlice_l173_71_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_71_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_71_3 = {1'd0, _zz_when_ArraySlice_l112_71};
  assign _zz_when_ArraySlice_l118_71_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_71 = _zz_when_ArraySlice_l118_71_1[5:0];
  assign _zz_when_ArraySlice_l173_71_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_71_1 = {3'd0, _zz_when_ArraySlice_l173_71_2};
  assign _zz_when_ArraySlice_l173_71_3 = (_zz_when_ArraySlice_l173_71_4 + _zz_when_ArraySlice_l173_71_8);
  assign _zz_when_ArraySlice_l173_71_4 = (_zz_when_ArraySlice_l173_71 - _zz_when_ArraySlice_l173_71_5);
  assign _zz_when_ArraySlice_l173_71_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_71_7);
  assign _zz_when_ArraySlice_l173_71_5 = {1'd0, _zz_when_ArraySlice_l173_71_6};
  assign _zz_when_ArraySlice_l173_71_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_71_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l421_2_1 = (_zz_when_ArraySlice_l421_2_2 + _zz_when_ArraySlice_l421_2_7);
  assign _zz_when_ArraySlice_l421_2_2 = (_zz_when_ArraySlice_l421_2_3 + _zz_when_ArraySlice_l421_2_5);
  assign _zz_when_ArraySlice_l421_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l421_2_4);
  assign _zz_when_ArraySlice_l421_2_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l421_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l421_2_5 = {5'd0, _zz_when_ArraySlice_l421_2_6};
  assign _zz_when_ArraySlice_l421_2_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l421_2_7 = {1'd0, _zz_when_ArraySlice_l421_2_8};
  assign _zz_selectReadFifo_2_25 = 1'b1;
  assign _zz_selectReadFifo_2_24 = {5'd0, _zz_selectReadFifo_2_25};
  assign _zz_when_ArraySlice_l425_2_1 = (_zz_when_ArraySlice_l425_2_2 % aReg);
  assign _zz_when_ArraySlice_l425_2_2 = (handshakeTimes_2_value + _zz_when_ArraySlice_l425_2_3);
  assign _zz_when_ArraySlice_l425_2_4 = 1'b1;
  assign _zz_when_ArraySlice_l425_2_3 = {12'd0, _zz_when_ArraySlice_l425_2_4};
  assign _zz_when_ArraySlice_l436_2_2 = (_zz_when_ArraySlice_l436_2_3 - _zz_when_ArraySlice_l436_2_4);
  assign _zz_when_ArraySlice_l436_2_1 = {7'd0, _zz_when_ArraySlice_l436_2_2};
  assign _zz_when_ArraySlice_l436_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l436_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l436_2_4 = {5'd0, _zz_when_ArraySlice_l436_2_5};
  assign _zz__zz_when_ArraySlice_l94_8 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_8 = (_zz_when_ArraySlice_l95_8_1 - _zz_when_ArraySlice_l95_8_4);
  assign _zz_when_ArraySlice_l95_8_1 = (_zz_when_ArraySlice_l95_8_2 + _zz_when_ArraySlice_l95_8_3);
  assign _zz_when_ArraySlice_l95_8_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_8_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_8_4 = {1'd0, _zz_when_ArraySlice_l94_8};
  assign _zz__zz_when_ArraySlice_l437_2_1 = (_zz__zz_when_ArraySlice_l437_2_2 + _zz__zz_when_ArraySlice_l437_2_3);
  assign _zz__zz_when_ArraySlice_l437_2_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l437_2_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l437_2_4 = {1'd0, _zz_when_ArraySlice_l94_8};
  assign _zz_when_ArraySlice_l99_8_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_8 = _zz_when_ArraySlice_l99_8_1[5:0];
  assign _zz_when_ArraySlice_l437_2_1 = (outSliceNumb_2_value + _zz_when_ArraySlice_l437_2_2);
  assign _zz_when_ArraySlice_l437_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l437_2_2 = {6'd0, _zz_when_ArraySlice_l437_2_3};
  assign _zz_when_ArraySlice_l437_2_4 = (_zz_when_ArraySlice_l437_2 / aReg);
  assign _zz_selectReadFifo_2_26 = (selectReadFifo_2 - _zz_selectReadFifo_2_27);
  assign _zz_selectReadFifo_2_27 = {3'd0, bReg};
  assign _zz_selectReadFifo_2_29 = 1'b1;
  assign _zz_selectReadFifo_2_28 = {5'd0, _zz_selectReadFifo_2_29};
  assign _zz_when_ArraySlice_l165_72 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_72_1);
  assign _zz_when_ArraySlice_l165_72_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_72_1 = {3'd0, _zz_when_ArraySlice_l165_72_2};
  assign _zz_when_ArraySlice_l166_72 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_72_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_72_3);
  assign _zz_when_ArraySlice_l166_72_1 = {1'd0, _zz_when_ArraySlice_l166_72_2};
  assign _zz_when_ArraySlice_l166_72_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_72_4);
  assign _zz_when_ArraySlice_l166_72_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_72_4 = {3'd0, _zz_when_ArraySlice_l166_72_5};
  assign _zz__zz_when_ArraySlice_l112_72 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_72 = (_zz_when_ArraySlice_l113_72_1 - _zz_when_ArraySlice_l113_72_4);
  assign _zz_when_ArraySlice_l113_72_1 = (_zz_when_ArraySlice_l113_72_2 + _zz_when_ArraySlice_l113_72_3);
  assign _zz_when_ArraySlice_l113_72_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_72_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_72_4 = {1'd0, _zz_when_ArraySlice_l112_72};
  assign _zz__zz_when_ArraySlice_l173_72 = (_zz__zz_when_ArraySlice_l173_72_1 + _zz__zz_when_ArraySlice_l173_72_2);
  assign _zz__zz_when_ArraySlice_l173_72_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_72_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_72_3 = {1'd0, _zz_when_ArraySlice_l112_72};
  assign _zz_when_ArraySlice_l118_72_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_72 = _zz_when_ArraySlice_l118_72_1[5:0];
  assign _zz_when_ArraySlice_l173_72_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_72_2 = (_zz_when_ArraySlice_l173_72_3 + _zz_when_ArraySlice_l173_72_8);
  assign _zz_when_ArraySlice_l173_72_3 = (_zz_when_ArraySlice_l173_72 - _zz_when_ArraySlice_l173_72_4);
  assign _zz_when_ArraySlice_l173_72_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_72_6);
  assign _zz_when_ArraySlice_l173_72_4 = {1'd0, _zz_when_ArraySlice_l173_72_5};
  assign _zz_when_ArraySlice_l173_72_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_72_6 = {3'd0, _zz_when_ArraySlice_l173_72_7};
  assign _zz_when_ArraySlice_l173_72_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_73 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_73_1);
  assign _zz_when_ArraySlice_l165_73_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_73_1 = {2'd0, _zz_when_ArraySlice_l165_73_2};
  assign _zz_when_ArraySlice_l166_73 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_73_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_73_2);
  assign _zz_when_ArraySlice_l166_73_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_73_3);
  assign _zz_when_ArraySlice_l166_73_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_73_3 = {2'd0, _zz_when_ArraySlice_l166_73_4};
  assign _zz__zz_when_ArraySlice_l112_73 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_73 = (_zz_when_ArraySlice_l113_73_1 - _zz_when_ArraySlice_l113_73_4);
  assign _zz_when_ArraySlice_l113_73_1 = (_zz_when_ArraySlice_l113_73_2 + _zz_when_ArraySlice_l113_73_3);
  assign _zz_when_ArraySlice_l113_73_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_73_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_73_4 = {1'd0, _zz_when_ArraySlice_l112_73};
  assign _zz__zz_when_ArraySlice_l173_73 = (_zz__zz_when_ArraySlice_l173_73_1 + _zz__zz_when_ArraySlice_l173_73_2);
  assign _zz__zz_when_ArraySlice_l173_73_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_73_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_73_3 = {1'd0, _zz_when_ArraySlice_l112_73};
  assign _zz_when_ArraySlice_l118_73_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_73 = _zz_when_ArraySlice_l118_73_1[5:0];
  assign _zz_when_ArraySlice_l173_73_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_73_1 = {1'd0, _zz_when_ArraySlice_l173_73_2};
  assign _zz_when_ArraySlice_l173_73_3 = (_zz_when_ArraySlice_l173_73_4 + _zz_when_ArraySlice_l173_73_9);
  assign _zz_when_ArraySlice_l173_73_4 = (_zz_when_ArraySlice_l173_73 - _zz_when_ArraySlice_l173_73_5);
  assign _zz_when_ArraySlice_l173_73_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_73_7);
  assign _zz_when_ArraySlice_l173_73_5 = {1'd0, _zz_when_ArraySlice_l173_73_6};
  assign _zz_when_ArraySlice_l173_73_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_73_7 = {2'd0, _zz_when_ArraySlice_l173_73_8};
  assign _zz_when_ArraySlice_l173_73_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_74 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_74_1);
  assign _zz_when_ArraySlice_l165_74_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_74_1 = {1'd0, _zz_when_ArraySlice_l165_74_2};
  assign _zz_when_ArraySlice_l166_74 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_74_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_74_2);
  assign _zz_when_ArraySlice_l166_74_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_74_3);
  assign _zz_when_ArraySlice_l166_74_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_74_3 = {1'd0, _zz_when_ArraySlice_l166_74_4};
  assign _zz__zz_when_ArraySlice_l112_74 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_74 = (_zz_when_ArraySlice_l113_74_1 - _zz_when_ArraySlice_l113_74_4);
  assign _zz_when_ArraySlice_l113_74_1 = (_zz_when_ArraySlice_l113_74_2 + _zz_when_ArraySlice_l113_74_3);
  assign _zz_when_ArraySlice_l113_74_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_74_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_74_4 = {1'd0, _zz_when_ArraySlice_l112_74};
  assign _zz__zz_when_ArraySlice_l173_74 = (_zz__zz_when_ArraySlice_l173_74_1 + _zz__zz_when_ArraySlice_l173_74_2);
  assign _zz__zz_when_ArraySlice_l173_74_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_74_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_74_3 = {1'd0, _zz_when_ArraySlice_l112_74};
  assign _zz_when_ArraySlice_l118_74_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_74 = _zz_when_ArraySlice_l118_74_1[5:0];
  assign _zz_when_ArraySlice_l173_74_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_74_1 = {1'd0, _zz_when_ArraySlice_l173_74_2};
  assign _zz_when_ArraySlice_l173_74_3 = (_zz_when_ArraySlice_l173_74_4 + _zz_when_ArraySlice_l173_74_9);
  assign _zz_when_ArraySlice_l173_74_4 = (_zz_when_ArraySlice_l173_74 - _zz_when_ArraySlice_l173_74_5);
  assign _zz_when_ArraySlice_l173_74_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_74_7);
  assign _zz_when_ArraySlice_l173_74_5 = {1'd0, _zz_when_ArraySlice_l173_74_6};
  assign _zz_when_ArraySlice_l173_74_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_74_7 = {1'd0, _zz_when_ArraySlice_l173_74_8};
  assign _zz_when_ArraySlice_l173_74_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_75 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_75_1);
  assign _zz_when_ArraySlice_l165_75_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_75_1 = {1'd0, _zz_when_ArraySlice_l165_75_2};
  assign _zz_when_ArraySlice_l166_75 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_75_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_75_2);
  assign _zz_when_ArraySlice_l166_75_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_75_3);
  assign _zz_when_ArraySlice_l166_75_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_75_3 = {1'd0, _zz_when_ArraySlice_l166_75_4};
  assign _zz__zz_when_ArraySlice_l112_75 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_75 = (_zz_when_ArraySlice_l113_75_1 - _zz_when_ArraySlice_l113_75_4);
  assign _zz_when_ArraySlice_l113_75_1 = (_zz_when_ArraySlice_l113_75_2 + _zz_when_ArraySlice_l113_75_3);
  assign _zz_when_ArraySlice_l113_75_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_75_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_75_4 = {1'd0, _zz_when_ArraySlice_l112_75};
  assign _zz__zz_when_ArraySlice_l173_75 = (_zz__zz_when_ArraySlice_l173_75_1 + _zz__zz_when_ArraySlice_l173_75_2);
  assign _zz__zz_when_ArraySlice_l173_75_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_75_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_75_3 = {1'd0, _zz_when_ArraySlice_l112_75};
  assign _zz_when_ArraySlice_l118_75_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_75 = _zz_when_ArraySlice_l118_75_1[5:0];
  assign _zz_when_ArraySlice_l173_75_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_75_1 = {1'd0, _zz_when_ArraySlice_l173_75_2};
  assign _zz_when_ArraySlice_l173_75_3 = (_zz_when_ArraySlice_l173_75_4 + _zz_when_ArraySlice_l173_75_9);
  assign _zz_when_ArraySlice_l173_75_4 = (_zz_when_ArraySlice_l173_75 - _zz_when_ArraySlice_l173_75_5);
  assign _zz_when_ArraySlice_l173_75_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_75_7);
  assign _zz_when_ArraySlice_l173_75_5 = {1'd0, _zz_when_ArraySlice_l173_75_6};
  assign _zz_when_ArraySlice_l173_75_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_75_7 = {1'd0, _zz_when_ArraySlice_l173_75_8};
  assign _zz_when_ArraySlice_l173_75_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_76 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_76_1);
  assign _zz_when_ArraySlice_l165_76_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_76 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_76_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_76_2);
  assign _zz_when_ArraySlice_l166_76_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_76_3);
  assign _zz_when_ArraySlice_l166_76_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_76 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_76 = (_zz_when_ArraySlice_l113_76_1 - _zz_when_ArraySlice_l113_76_4);
  assign _zz_when_ArraySlice_l113_76_1 = (_zz_when_ArraySlice_l113_76_2 + _zz_when_ArraySlice_l113_76_3);
  assign _zz_when_ArraySlice_l113_76_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_76_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_76_4 = {1'd0, _zz_when_ArraySlice_l112_76};
  assign _zz__zz_when_ArraySlice_l173_76 = (_zz__zz_when_ArraySlice_l173_76_1 + _zz__zz_when_ArraySlice_l173_76_2);
  assign _zz__zz_when_ArraySlice_l173_76_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_76_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_76_3 = {1'd0, _zz_when_ArraySlice_l112_76};
  assign _zz_when_ArraySlice_l118_76_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_76 = _zz_when_ArraySlice_l118_76_1[5:0];
  assign _zz_when_ArraySlice_l173_76_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_76_1 = {1'd0, _zz_when_ArraySlice_l173_76_2};
  assign _zz_when_ArraySlice_l173_76_3 = (_zz_when_ArraySlice_l173_76_4 + _zz_when_ArraySlice_l173_76_8);
  assign _zz_when_ArraySlice_l173_76_4 = (_zz_when_ArraySlice_l173_76 - _zz_when_ArraySlice_l173_76_5);
  assign _zz_when_ArraySlice_l173_76_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_76_7);
  assign _zz_when_ArraySlice_l173_76_5 = {1'd0, _zz_when_ArraySlice_l173_76_6};
  assign _zz_when_ArraySlice_l173_76_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_76_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_77 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_77_1);
  assign _zz_when_ArraySlice_l165_77_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_77_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_77 = {1'd0, _zz_when_ArraySlice_l166_77_1};
  assign _zz_when_ArraySlice_l166_77_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_77_3);
  assign _zz_when_ArraySlice_l166_77_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_77_4);
  assign _zz_when_ArraySlice_l166_77_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_77 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_77 = (_zz_when_ArraySlice_l113_77_1 - _zz_when_ArraySlice_l113_77_4);
  assign _zz_when_ArraySlice_l113_77_1 = (_zz_when_ArraySlice_l113_77_2 + _zz_when_ArraySlice_l113_77_3);
  assign _zz_when_ArraySlice_l113_77_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_77_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_77_4 = {1'd0, _zz_when_ArraySlice_l112_77};
  assign _zz__zz_when_ArraySlice_l173_77 = (_zz__zz_when_ArraySlice_l173_77_1 + _zz__zz_when_ArraySlice_l173_77_2);
  assign _zz__zz_when_ArraySlice_l173_77_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_77_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_77_3 = {1'd0, _zz_when_ArraySlice_l112_77};
  assign _zz_when_ArraySlice_l118_77_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_77 = _zz_when_ArraySlice_l118_77_1[5:0];
  assign _zz_when_ArraySlice_l173_77_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_77_1 = {2'd0, _zz_when_ArraySlice_l173_77_2};
  assign _zz_when_ArraySlice_l173_77_3 = (_zz_when_ArraySlice_l173_77_4 + _zz_when_ArraySlice_l173_77_8);
  assign _zz_when_ArraySlice_l173_77_4 = (_zz_when_ArraySlice_l173_77 - _zz_when_ArraySlice_l173_77_5);
  assign _zz_when_ArraySlice_l173_77_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_77_7);
  assign _zz_when_ArraySlice_l173_77_5 = {1'd0, _zz_when_ArraySlice_l173_77_6};
  assign _zz_when_ArraySlice_l173_77_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_77_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_78 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_78_1);
  assign _zz_when_ArraySlice_l165_78_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_78_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_78 = {1'd0, _zz_when_ArraySlice_l166_78_1};
  assign _zz_when_ArraySlice_l166_78_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_78_3);
  assign _zz_when_ArraySlice_l166_78_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_78_4);
  assign _zz_when_ArraySlice_l166_78_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_78 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_78 = (_zz_when_ArraySlice_l113_78_1 - _zz_when_ArraySlice_l113_78_4);
  assign _zz_when_ArraySlice_l113_78_1 = (_zz_when_ArraySlice_l113_78_2 + _zz_when_ArraySlice_l113_78_3);
  assign _zz_when_ArraySlice_l113_78_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_78_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_78_4 = {1'd0, _zz_when_ArraySlice_l112_78};
  assign _zz__zz_when_ArraySlice_l173_78 = (_zz__zz_when_ArraySlice_l173_78_1 + _zz__zz_when_ArraySlice_l173_78_2);
  assign _zz__zz_when_ArraySlice_l173_78_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_78_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_78_3 = {1'd0, _zz_when_ArraySlice_l112_78};
  assign _zz_when_ArraySlice_l118_78_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_78 = _zz_when_ArraySlice_l118_78_1[5:0];
  assign _zz_when_ArraySlice_l173_78_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_78_1 = {2'd0, _zz_when_ArraySlice_l173_78_2};
  assign _zz_when_ArraySlice_l173_78_3 = (_zz_when_ArraySlice_l173_78_4 + _zz_when_ArraySlice_l173_78_8);
  assign _zz_when_ArraySlice_l173_78_4 = (_zz_when_ArraySlice_l173_78 - _zz_when_ArraySlice_l173_78_5);
  assign _zz_when_ArraySlice_l173_78_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_78_7);
  assign _zz_when_ArraySlice_l173_78_5 = {1'd0, _zz_when_ArraySlice_l173_78_6};
  assign _zz_when_ArraySlice_l173_78_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_78_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_79 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_79_1);
  assign _zz_when_ArraySlice_l165_79_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_79_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_79 = {2'd0, _zz_when_ArraySlice_l166_79_1};
  assign _zz_when_ArraySlice_l166_79_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_79_3);
  assign _zz_when_ArraySlice_l166_79_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_79_4);
  assign _zz_when_ArraySlice_l166_79_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_79 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_79 = (_zz_when_ArraySlice_l113_79_1 - _zz_when_ArraySlice_l113_79_4);
  assign _zz_when_ArraySlice_l113_79_1 = (_zz_when_ArraySlice_l113_79_2 + _zz_when_ArraySlice_l113_79_3);
  assign _zz_when_ArraySlice_l113_79_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_79_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_79_4 = {1'd0, _zz_when_ArraySlice_l112_79};
  assign _zz__zz_when_ArraySlice_l173_79 = (_zz__zz_when_ArraySlice_l173_79_1 + _zz__zz_when_ArraySlice_l173_79_2);
  assign _zz__zz_when_ArraySlice_l173_79_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_79_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_79_3 = {1'd0, _zz_when_ArraySlice_l112_79};
  assign _zz_when_ArraySlice_l118_79_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_79 = _zz_when_ArraySlice_l118_79_1[5:0];
  assign _zz_when_ArraySlice_l173_79_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_79_1 = {3'd0, _zz_when_ArraySlice_l173_79_2};
  assign _zz_when_ArraySlice_l173_79_3 = (_zz_when_ArraySlice_l173_79_4 + _zz_when_ArraySlice_l173_79_8);
  assign _zz_when_ArraySlice_l173_79_4 = (_zz_when_ArraySlice_l173_79 - _zz_when_ArraySlice_l173_79_5);
  assign _zz_when_ArraySlice_l173_79_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_79_7);
  assign _zz_when_ArraySlice_l173_79_5 = {1'd0, _zz_when_ArraySlice_l173_79_6};
  assign _zz_when_ArraySlice_l173_79_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_79_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_2_31 = 1'b1;
  assign _zz_selectReadFifo_2_30 = {5'd0, _zz_selectReadFifo_2_31};
  assign _zz_when_ArraySlice_l448_2_1 = (_zz_when_ArraySlice_l448_2_2 % aReg);
  assign _zz_when_ArraySlice_l448_2_2 = (handshakeTimes_2_value + _zz_when_ArraySlice_l448_2_3);
  assign _zz_when_ArraySlice_l448_2_4 = 1'b1;
  assign _zz_when_ArraySlice_l448_2_3 = {12'd0, _zz_when_ArraySlice_l448_2_4};
  assign _zz_when_ArraySlice_l434_2_1 = (selectReadFifo_2 + _zz_when_ArraySlice_l434_2_2);
  assign _zz_when_ArraySlice_l434_2_3 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l434_2_2 = {1'd0, _zz_when_ArraySlice_l434_2_3};
  assign _zz_when_ArraySlice_l455_2_2 = (_zz_when_ArraySlice_l455_2_3 - _zz_when_ArraySlice_l455_2_4);
  assign _zz_when_ArraySlice_l455_2_1 = {7'd0, _zz_when_ArraySlice_l455_2_2};
  assign _zz_when_ArraySlice_l455_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l455_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l455_2_4 = {5'd0, _zz_when_ArraySlice_l455_2_5};
  assign _zz_when_ArraySlice_l373_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l373_3_1);
  assign _zz_when_ArraySlice_l373_3_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l373_3_1 = {1'd0, _zz_when_ArraySlice_l373_3_2};
  assign _zz_when_ArraySlice_l374_3_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l374_3_3);
  assign _zz_when_ArraySlice_l374_3_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l374_3_3 = {1'd0, _zz_when_ArraySlice_l374_3_4};
  assign _zz__zz_outputStreamArrayData_3_valid_1 = (bReg * 2'b11);
  assign _zz__zz_outputStreamArrayData_3_valid = {1'd0, _zz__zz_outputStreamArrayData_3_valid_1};
  assign _zz_when_ArraySlice_l380_3_2 = 1'b1;
  assign _zz_when_ArraySlice_l380_3_1 = {6'd0, _zz_when_ArraySlice_l380_3_2};
  assign _zz_when_ArraySlice_l380_3_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l380_3_5);
  assign _zz_when_ArraySlice_l380_3_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l380_3_5 = {1'd0, _zz_when_ArraySlice_l380_3_6};
  assign _zz_when_ArraySlice_l381_3_2 = (_zz_when_ArraySlice_l381_3_3 - _zz_when_ArraySlice_l381_3_4);
  assign _zz_when_ArraySlice_l381_3_1 = {7'd0, _zz_when_ArraySlice_l381_3_2};
  assign _zz_when_ArraySlice_l381_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l381_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l381_3_4 = {5'd0, _zz_when_ArraySlice_l381_3_5};
  assign _zz_selectReadFifo_3 = (selectReadFifo_3 - _zz_selectReadFifo_3_1);
  assign _zz_selectReadFifo_3_1 = {3'd0, bReg};
  assign _zz_selectReadFifo_3_3 = 1'b1;
  assign _zz_selectReadFifo_3_2 = {5'd0, _zz_selectReadFifo_3_3};
  assign _zz_selectReadFifo_3_5 = 1'b1;
  assign _zz_selectReadFifo_3_4 = {5'd0, _zz_selectReadFifo_3_5};
  assign _zz_when_ArraySlice_l384_3_1 = (_zz_when_ArraySlice_l384_3_2 % aReg);
  assign _zz_when_ArraySlice_l384_3_2 = (handshakeTimes_3_value + _zz_when_ArraySlice_l384_3_3);
  assign _zz_when_ArraySlice_l384_3_4 = 1'b1;
  assign _zz_when_ArraySlice_l384_3_3 = {12'd0, _zz_when_ArraySlice_l384_3_4};
  assign _zz_when_ArraySlice_l389_3_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l389_3_3);
  assign _zz_when_ArraySlice_l389_3_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l389_3_3 = {1'd0, _zz_when_ArraySlice_l389_3_4};
  assign _zz_when_ArraySlice_l389_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l389_3_5 = {6'd0, _zz_when_ArraySlice_l389_3_6};
  assign _zz_when_ArraySlice_l390_3_2 = (_zz_when_ArraySlice_l390_3_3 - _zz_when_ArraySlice_l390_3_4);
  assign _zz_when_ArraySlice_l390_3_1 = {7'd0, _zz_when_ArraySlice_l390_3_2};
  assign _zz_when_ArraySlice_l390_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l390_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l390_3_4 = {5'd0, _zz_when_ArraySlice_l390_3_5};
  assign _zz__zz_when_ArraySlice_l94_9 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_9 = (_zz_when_ArraySlice_l95_9_1 - _zz_when_ArraySlice_l95_9_4);
  assign _zz_when_ArraySlice_l95_9_1 = (_zz_when_ArraySlice_l95_9_2 + _zz_when_ArraySlice_l95_9_3);
  assign _zz_when_ArraySlice_l95_9_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_9_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_9_4 = {1'd0, _zz_when_ArraySlice_l94_9};
  assign _zz__zz_when_ArraySlice_l392_3_1 = (_zz__zz_when_ArraySlice_l392_3_2 + _zz__zz_when_ArraySlice_l392_3_3);
  assign _zz__zz_when_ArraySlice_l392_3_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l392_3_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l392_3_4 = {1'd0, _zz_when_ArraySlice_l94_9};
  assign _zz_when_ArraySlice_l99_9_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_9 = _zz_when_ArraySlice_l99_9_1[5:0];
  assign _zz_when_ArraySlice_l392_3_1 = (outSliceNumb_3_value + _zz_when_ArraySlice_l392_3_2);
  assign _zz_when_ArraySlice_l392_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l392_3_2 = {6'd0, _zz_when_ArraySlice_l392_3_3};
  assign _zz_when_ArraySlice_l392_3_4 = (_zz_when_ArraySlice_l392_3 / aReg);
  assign _zz_selectReadFifo_3_6 = (selectReadFifo_3 - _zz_selectReadFifo_3_7);
  assign _zz_selectReadFifo_3_7 = {3'd0, bReg};
  assign _zz_selectReadFifo_3_9 = 1'b1;
  assign _zz_selectReadFifo_3_8 = {5'd0, _zz_selectReadFifo_3_9};
  assign _zz_selectReadFifo_3_10 = (selectReadFifo_3 + _zz_selectReadFifo_3_11);
  assign _zz_selectReadFifo_3_11 = (3'b111 * bReg);
  assign _zz_selectReadFifo_3_13 = 1'b1;
  assign _zz_selectReadFifo_3_12 = {5'd0, _zz_selectReadFifo_3_13};
  assign _zz_when_ArraySlice_l165_80 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_80_1);
  assign _zz_when_ArraySlice_l165_80_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_80_1 = {3'd0, _zz_when_ArraySlice_l165_80_2};
  assign _zz_when_ArraySlice_l166_80 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_80_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_80_3);
  assign _zz_when_ArraySlice_l166_80_1 = {1'd0, _zz_when_ArraySlice_l166_80_2};
  assign _zz_when_ArraySlice_l166_80_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_80_4);
  assign _zz_when_ArraySlice_l166_80_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_80_4 = {3'd0, _zz_when_ArraySlice_l166_80_5};
  assign _zz__zz_when_ArraySlice_l112_80 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_80 = (_zz_when_ArraySlice_l113_80_1 - _zz_when_ArraySlice_l113_80_4);
  assign _zz_when_ArraySlice_l113_80_1 = (_zz_when_ArraySlice_l113_80_2 + _zz_when_ArraySlice_l113_80_3);
  assign _zz_when_ArraySlice_l113_80_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_80_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_80_4 = {1'd0, _zz_when_ArraySlice_l112_80};
  assign _zz__zz_when_ArraySlice_l173_80 = (_zz__zz_when_ArraySlice_l173_80_1 + _zz__zz_when_ArraySlice_l173_80_2);
  assign _zz__zz_when_ArraySlice_l173_80_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_80_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_80_3 = {1'd0, _zz_when_ArraySlice_l112_80};
  assign _zz_when_ArraySlice_l118_80_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_80 = _zz_when_ArraySlice_l118_80_1[5:0];
  assign _zz_when_ArraySlice_l173_80_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_80_2 = (_zz_when_ArraySlice_l173_80_3 + _zz_when_ArraySlice_l173_80_8);
  assign _zz_when_ArraySlice_l173_80_3 = (_zz_when_ArraySlice_l173_80 - _zz_when_ArraySlice_l173_80_4);
  assign _zz_when_ArraySlice_l173_80_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_80_6);
  assign _zz_when_ArraySlice_l173_80_4 = {1'd0, _zz_when_ArraySlice_l173_80_5};
  assign _zz_when_ArraySlice_l173_80_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_80_6 = {3'd0, _zz_when_ArraySlice_l173_80_7};
  assign _zz_when_ArraySlice_l173_80_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_81 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_81_1);
  assign _zz_when_ArraySlice_l165_81_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_81_1 = {2'd0, _zz_when_ArraySlice_l165_81_2};
  assign _zz_when_ArraySlice_l166_81 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_81_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_81_2);
  assign _zz_when_ArraySlice_l166_81_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_81_3);
  assign _zz_when_ArraySlice_l166_81_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_81_3 = {2'd0, _zz_when_ArraySlice_l166_81_4};
  assign _zz__zz_when_ArraySlice_l112_81 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_81 = (_zz_when_ArraySlice_l113_81_1 - _zz_when_ArraySlice_l113_81_4);
  assign _zz_when_ArraySlice_l113_81_1 = (_zz_when_ArraySlice_l113_81_2 + _zz_when_ArraySlice_l113_81_3);
  assign _zz_when_ArraySlice_l113_81_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_81_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_81_4 = {1'd0, _zz_when_ArraySlice_l112_81};
  assign _zz__zz_when_ArraySlice_l173_81 = (_zz__zz_when_ArraySlice_l173_81_1 + _zz__zz_when_ArraySlice_l173_81_2);
  assign _zz__zz_when_ArraySlice_l173_81_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_81_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_81_3 = {1'd0, _zz_when_ArraySlice_l112_81};
  assign _zz_when_ArraySlice_l118_81_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_81 = _zz_when_ArraySlice_l118_81_1[5:0];
  assign _zz_when_ArraySlice_l173_81_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_81_1 = {1'd0, _zz_when_ArraySlice_l173_81_2};
  assign _zz_when_ArraySlice_l173_81_3 = (_zz_when_ArraySlice_l173_81_4 + _zz_when_ArraySlice_l173_81_9);
  assign _zz_when_ArraySlice_l173_81_4 = (_zz_when_ArraySlice_l173_81 - _zz_when_ArraySlice_l173_81_5);
  assign _zz_when_ArraySlice_l173_81_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_81_7);
  assign _zz_when_ArraySlice_l173_81_5 = {1'd0, _zz_when_ArraySlice_l173_81_6};
  assign _zz_when_ArraySlice_l173_81_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_81_7 = {2'd0, _zz_when_ArraySlice_l173_81_8};
  assign _zz_when_ArraySlice_l173_81_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_82 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_82_1);
  assign _zz_when_ArraySlice_l165_82_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_82_1 = {1'd0, _zz_when_ArraySlice_l165_82_2};
  assign _zz_when_ArraySlice_l166_82 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_82_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_82_2);
  assign _zz_when_ArraySlice_l166_82_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_82_3);
  assign _zz_when_ArraySlice_l166_82_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_82_3 = {1'd0, _zz_when_ArraySlice_l166_82_4};
  assign _zz__zz_when_ArraySlice_l112_82 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_82 = (_zz_when_ArraySlice_l113_82_1 - _zz_when_ArraySlice_l113_82_4);
  assign _zz_when_ArraySlice_l113_82_1 = (_zz_when_ArraySlice_l113_82_2 + _zz_when_ArraySlice_l113_82_3);
  assign _zz_when_ArraySlice_l113_82_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_82_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_82_4 = {1'd0, _zz_when_ArraySlice_l112_82};
  assign _zz__zz_when_ArraySlice_l173_82 = (_zz__zz_when_ArraySlice_l173_82_1 + _zz__zz_when_ArraySlice_l173_82_2);
  assign _zz__zz_when_ArraySlice_l173_82_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_82_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_82_3 = {1'd0, _zz_when_ArraySlice_l112_82};
  assign _zz_when_ArraySlice_l118_82_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_82 = _zz_when_ArraySlice_l118_82_1[5:0];
  assign _zz_when_ArraySlice_l173_82_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_82_1 = {1'd0, _zz_when_ArraySlice_l173_82_2};
  assign _zz_when_ArraySlice_l173_82_3 = (_zz_when_ArraySlice_l173_82_4 + _zz_when_ArraySlice_l173_82_9);
  assign _zz_when_ArraySlice_l173_82_4 = (_zz_when_ArraySlice_l173_82 - _zz_when_ArraySlice_l173_82_5);
  assign _zz_when_ArraySlice_l173_82_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_82_7);
  assign _zz_when_ArraySlice_l173_82_5 = {1'd0, _zz_when_ArraySlice_l173_82_6};
  assign _zz_when_ArraySlice_l173_82_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_82_7 = {1'd0, _zz_when_ArraySlice_l173_82_8};
  assign _zz_when_ArraySlice_l173_82_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_83 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_83_1);
  assign _zz_when_ArraySlice_l165_83_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_83_1 = {1'd0, _zz_when_ArraySlice_l165_83_2};
  assign _zz_when_ArraySlice_l166_83 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_83_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_83_2);
  assign _zz_when_ArraySlice_l166_83_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_83_3);
  assign _zz_when_ArraySlice_l166_83_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_83_3 = {1'd0, _zz_when_ArraySlice_l166_83_4};
  assign _zz__zz_when_ArraySlice_l112_83 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_83 = (_zz_when_ArraySlice_l113_83_1 - _zz_when_ArraySlice_l113_83_4);
  assign _zz_when_ArraySlice_l113_83_1 = (_zz_when_ArraySlice_l113_83_2 + _zz_when_ArraySlice_l113_83_3);
  assign _zz_when_ArraySlice_l113_83_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_83_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_83_4 = {1'd0, _zz_when_ArraySlice_l112_83};
  assign _zz__zz_when_ArraySlice_l173_83 = (_zz__zz_when_ArraySlice_l173_83_1 + _zz__zz_when_ArraySlice_l173_83_2);
  assign _zz__zz_when_ArraySlice_l173_83_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_83_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_83_3 = {1'd0, _zz_when_ArraySlice_l112_83};
  assign _zz_when_ArraySlice_l118_83_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_83 = _zz_when_ArraySlice_l118_83_1[5:0];
  assign _zz_when_ArraySlice_l173_83_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_83_1 = {1'd0, _zz_when_ArraySlice_l173_83_2};
  assign _zz_when_ArraySlice_l173_83_3 = (_zz_when_ArraySlice_l173_83_4 + _zz_when_ArraySlice_l173_83_9);
  assign _zz_when_ArraySlice_l173_83_4 = (_zz_when_ArraySlice_l173_83 - _zz_when_ArraySlice_l173_83_5);
  assign _zz_when_ArraySlice_l173_83_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_83_7);
  assign _zz_when_ArraySlice_l173_83_5 = {1'd0, _zz_when_ArraySlice_l173_83_6};
  assign _zz_when_ArraySlice_l173_83_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_83_7 = {1'd0, _zz_when_ArraySlice_l173_83_8};
  assign _zz_when_ArraySlice_l173_83_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_84 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_84_1);
  assign _zz_when_ArraySlice_l165_84_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_84 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_84_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_84_2);
  assign _zz_when_ArraySlice_l166_84_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_84_3);
  assign _zz_when_ArraySlice_l166_84_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_84 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_84 = (_zz_when_ArraySlice_l113_84_1 - _zz_when_ArraySlice_l113_84_4);
  assign _zz_when_ArraySlice_l113_84_1 = (_zz_when_ArraySlice_l113_84_2 + _zz_when_ArraySlice_l113_84_3);
  assign _zz_when_ArraySlice_l113_84_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_84_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_84_4 = {1'd0, _zz_when_ArraySlice_l112_84};
  assign _zz__zz_when_ArraySlice_l173_84 = (_zz__zz_when_ArraySlice_l173_84_1 + _zz__zz_when_ArraySlice_l173_84_2);
  assign _zz__zz_when_ArraySlice_l173_84_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_84_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_84_3 = {1'd0, _zz_when_ArraySlice_l112_84};
  assign _zz_when_ArraySlice_l118_84_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_84 = _zz_when_ArraySlice_l118_84_1[5:0];
  assign _zz_when_ArraySlice_l173_84_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_84_1 = {1'd0, _zz_when_ArraySlice_l173_84_2};
  assign _zz_when_ArraySlice_l173_84_3 = (_zz_when_ArraySlice_l173_84_4 + _zz_when_ArraySlice_l173_84_8);
  assign _zz_when_ArraySlice_l173_84_4 = (_zz_when_ArraySlice_l173_84 - _zz_when_ArraySlice_l173_84_5);
  assign _zz_when_ArraySlice_l173_84_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_84_7);
  assign _zz_when_ArraySlice_l173_84_5 = {1'd0, _zz_when_ArraySlice_l173_84_6};
  assign _zz_when_ArraySlice_l173_84_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_84_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_85 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_85_1);
  assign _zz_when_ArraySlice_l165_85_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_85_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_85 = {1'd0, _zz_when_ArraySlice_l166_85_1};
  assign _zz_when_ArraySlice_l166_85_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_85_3);
  assign _zz_when_ArraySlice_l166_85_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_85_4);
  assign _zz_when_ArraySlice_l166_85_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_85 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_85 = (_zz_when_ArraySlice_l113_85_1 - _zz_when_ArraySlice_l113_85_4);
  assign _zz_when_ArraySlice_l113_85_1 = (_zz_when_ArraySlice_l113_85_2 + _zz_when_ArraySlice_l113_85_3);
  assign _zz_when_ArraySlice_l113_85_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_85_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_85_4 = {1'd0, _zz_when_ArraySlice_l112_85};
  assign _zz__zz_when_ArraySlice_l173_85 = (_zz__zz_when_ArraySlice_l173_85_1 + _zz__zz_when_ArraySlice_l173_85_2);
  assign _zz__zz_when_ArraySlice_l173_85_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_85_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_85_3 = {1'd0, _zz_when_ArraySlice_l112_85};
  assign _zz_when_ArraySlice_l118_85_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_85 = _zz_when_ArraySlice_l118_85_1[5:0];
  assign _zz_when_ArraySlice_l173_85_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_85_1 = {2'd0, _zz_when_ArraySlice_l173_85_2};
  assign _zz_when_ArraySlice_l173_85_3 = (_zz_when_ArraySlice_l173_85_4 + _zz_when_ArraySlice_l173_85_8);
  assign _zz_when_ArraySlice_l173_85_4 = (_zz_when_ArraySlice_l173_85 - _zz_when_ArraySlice_l173_85_5);
  assign _zz_when_ArraySlice_l173_85_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_85_7);
  assign _zz_when_ArraySlice_l173_85_5 = {1'd0, _zz_when_ArraySlice_l173_85_6};
  assign _zz_when_ArraySlice_l173_85_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_85_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_86 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_86_1);
  assign _zz_when_ArraySlice_l165_86_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_86_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_86 = {1'd0, _zz_when_ArraySlice_l166_86_1};
  assign _zz_when_ArraySlice_l166_86_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_86_3);
  assign _zz_when_ArraySlice_l166_86_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_86_4);
  assign _zz_when_ArraySlice_l166_86_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_86 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_86 = (_zz_when_ArraySlice_l113_86_1 - _zz_when_ArraySlice_l113_86_4);
  assign _zz_when_ArraySlice_l113_86_1 = (_zz_when_ArraySlice_l113_86_2 + _zz_when_ArraySlice_l113_86_3);
  assign _zz_when_ArraySlice_l113_86_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_86_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_86_4 = {1'd0, _zz_when_ArraySlice_l112_86};
  assign _zz__zz_when_ArraySlice_l173_86 = (_zz__zz_when_ArraySlice_l173_86_1 + _zz__zz_when_ArraySlice_l173_86_2);
  assign _zz__zz_when_ArraySlice_l173_86_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_86_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_86_3 = {1'd0, _zz_when_ArraySlice_l112_86};
  assign _zz_when_ArraySlice_l118_86_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_86 = _zz_when_ArraySlice_l118_86_1[5:0];
  assign _zz_when_ArraySlice_l173_86_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_86_1 = {2'd0, _zz_when_ArraySlice_l173_86_2};
  assign _zz_when_ArraySlice_l173_86_3 = (_zz_when_ArraySlice_l173_86_4 + _zz_when_ArraySlice_l173_86_8);
  assign _zz_when_ArraySlice_l173_86_4 = (_zz_when_ArraySlice_l173_86 - _zz_when_ArraySlice_l173_86_5);
  assign _zz_when_ArraySlice_l173_86_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_86_7);
  assign _zz_when_ArraySlice_l173_86_5 = {1'd0, _zz_when_ArraySlice_l173_86_6};
  assign _zz_when_ArraySlice_l173_86_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_86_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_87 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_87_1);
  assign _zz_when_ArraySlice_l165_87_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_87_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_87 = {2'd0, _zz_when_ArraySlice_l166_87_1};
  assign _zz_when_ArraySlice_l166_87_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_87_3);
  assign _zz_when_ArraySlice_l166_87_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_87_4);
  assign _zz_when_ArraySlice_l166_87_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_87 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_87 = (_zz_when_ArraySlice_l113_87_1 - _zz_when_ArraySlice_l113_87_4);
  assign _zz_when_ArraySlice_l113_87_1 = (_zz_when_ArraySlice_l113_87_2 + _zz_when_ArraySlice_l113_87_3);
  assign _zz_when_ArraySlice_l113_87_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_87_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_87_4 = {1'd0, _zz_when_ArraySlice_l112_87};
  assign _zz__zz_when_ArraySlice_l173_87 = (_zz__zz_when_ArraySlice_l173_87_1 + _zz__zz_when_ArraySlice_l173_87_2);
  assign _zz__zz_when_ArraySlice_l173_87_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_87_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_87_3 = {1'd0, _zz_when_ArraySlice_l112_87};
  assign _zz_when_ArraySlice_l118_87_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_87 = _zz_when_ArraySlice_l118_87_1[5:0];
  assign _zz_when_ArraySlice_l173_87_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_87_1 = {3'd0, _zz_when_ArraySlice_l173_87_2};
  assign _zz_when_ArraySlice_l173_87_3 = (_zz_when_ArraySlice_l173_87_4 + _zz_when_ArraySlice_l173_87_8);
  assign _zz_when_ArraySlice_l173_87_4 = (_zz_when_ArraySlice_l173_87 - _zz_when_ArraySlice_l173_87_5);
  assign _zz_when_ArraySlice_l173_87_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_87_7);
  assign _zz_when_ArraySlice_l173_87_5 = {1'd0, _zz_when_ArraySlice_l173_87_6};
  assign _zz_when_ArraySlice_l173_87_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_87_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l401_3_1 = (_zz_when_ArraySlice_l401_3_2 + _zz_when_ArraySlice_l401_3_7);
  assign _zz_when_ArraySlice_l401_3_2 = (_zz_when_ArraySlice_l401_3_3 + _zz_when_ArraySlice_l401_3_5);
  assign _zz_when_ArraySlice_l401_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l401_3_4);
  assign _zz_when_ArraySlice_l401_3_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l401_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l401_3_5 = {5'd0, _zz_when_ArraySlice_l401_3_6};
  assign _zz_when_ArraySlice_l401_3_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l401_3_7 = {1'd0, _zz_when_ArraySlice_l401_3_8};
  assign _zz_selectReadFifo_3_15 = 1'b1;
  assign _zz_selectReadFifo_3_14 = {5'd0, _zz_selectReadFifo_3_15};
  assign _zz_when_ArraySlice_l405_3_1 = (_zz_when_ArraySlice_l405_3_2 % aReg);
  assign _zz_when_ArraySlice_l405_3_2 = (handshakeTimes_3_value + _zz_when_ArraySlice_l405_3_3);
  assign _zz_when_ArraySlice_l405_3_4 = 1'b1;
  assign _zz_when_ArraySlice_l405_3_3 = {12'd0, _zz_when_ArraySlice_l405_3_4};
  assign _zz_when_ArraySlice_l409_3_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l409_3_3);
  assign _zz_when_ArraySlice_l409_3_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l409_3_3 = {1'd0, _zz_when_ArraySlice_l409_3_4};
  assign _zz_when_ArraySlice_l410_3_2 = (_zz_when_ArraySlice_l410_3_3 - _zz_when_ArraySlice_l410_3_4);
  assign _zz_when_ArraySlice_l410_3_1 = {7'd0, _zz_when_ArraySlice_l410_3_2};
  assign _zz_when_ArraySlice_l410_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l410_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l410_3_4 = {5'd0, _zz_when_ArraySlice_l410_3_5};
  assign _zz__zz_when_ArraySlice_l94_10 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_10 = (_zz_when_ArraySlice_l95_10_1 - _zz_when_ArraySlice_l95_10_4);
  assign _zz_when_ArraySlice_l95_10_1 = (_zz_when_ArraySlice_l95_10_2 + _zz_when_ArraySlice_l95_10_3);
  assign _zz_when_ArraySlice_l95_10_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_10_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_10_4 = {1'd0, _zz_when_ArraySlice_l94_10};
  assign _zz__zz_when_ArraySlice_l412_3_1 = (_zz__zz_when_ArraySlice_l412_3_2 + _zz__zz_when_ArraySlice_l412_3_3);
  assign _zz__zz_when_ArraySlice_l412_3_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l412_3_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l412_3_4 = {1'd0, _zz_when_ArraySlice_l94_10};
  assign _zz_when_ArraySlice_l99_10_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_10 = _zz_when_ArraySlice_l99_10_1[5:0];
  assign _zz_when_ArraySlice_l412_3_1 = (outSliceNumb_3_value + _zz_when_ArraySlice_l412_3_2);
  assign _zz_when_ArraySlice_l412_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l412_3_2 = {6'd0, _zz_when_ArraySlice_l412_3_3};
  assign _zz_when_ArraySlice_l412_3_4 = (_zz_when_ArraySlice_l412_3 / aReg);
  assign _zz_selectReadFifo_3_16 = (selectReadFifo_3 - _zz_selectReadFifo_3_17);
  assign _zz_selectReadFifo_3_17 = {3'd0, bReg};
  assign _zz_selectReadFifo_3_19 = 1'b1;
  assign _zz_selectReadFifo_3_18 = {5'd0, _zz_selectReadFifo_3_19};
  assign _zz_selectReadFifo_3_20 = (selectReadFifo_3 + _zz_selectReadFifo_3_21);
  assign _zz_selectReadFifo_3_21 = (3'b111 * bReg);
  assign _zz_selectReadFifo_3_23 = 1'b1;
  assign _zz_selectReadFifo_3_22 = {5'd0, _zz_selectReadFifo_3_23};
  assign _zz_when_ArraySlice_l165_88 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_88_1);
  assign _zz_when_ArraySlice_l165_88_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_88_1 = {3'd0, _zz_when_ArraySlice_l165_88_2};
  assign _zz_when_ArraySlice_l166_88 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_88_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_88_3);
  assign _zz_when_ArraySlice_l166_88_1 = {1'd0, _zz_when_ArraySlice_l166_88_2};
  assign _zz_when_ArraySlice_l166_88_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_88_4);
  assign _zz_when_ArraySlice_l166_88_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_88_4 = {3'd0, _zz_when_ArraySlice_l166_88_5};
  assign _zz__zz_when_ArraySlice_l112_88 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_88 = (_zz_when_ArraySlice_l113_88_1 - _zz_when_ArraySlice_l113_88_4);
  assign _zz_when_ArraySlice_l113_88_1 = (_zz_when_ArraySlice_l113_88_2 + _zz_when_ArraySlice_l113_88_3);
  assign _zz_when_ArraySlice_l113_88_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_88_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_88_4 = {1'd0, _zz_when_ArraySlice_l112_88};
  assign _zz__zz_when_ArraySlice_l173_88 = (_zz__zz_when_ArraySlice_l173_88_1 + _zz__zz_when_ArraySlice_l173_88_2);
  assign _zz__zz_when_ArraySlice_l173_88_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_88_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_88_3 = {1'd0, _zz_when_ArraySlice_l112_88};
  assign _zz_when_ArraySlice_l118_88_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_88 = _zz_when_ArraySlice_l118_88_1[5:0];
  assign _zz_when_ArraySlice_l173_88_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_88_2 = (_zz_when_ArraySlice_l173_88_3 + _zz_when_ArraySlice_l173_88_8);
  assign _zz_when_ArraySlice_l173_88_3 = (_zz_when_ArraySlice_l173_88 - _zz_when_ArraySlice_l173_88_4);
  assign _zz_when_ArraySlice_l173_88_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_88_6);
  assign _zz_when_ArraySlice_l173_88_4 = {1'd0, _zz_when_ArraySlice_l173_88_5};
  assign _zz_when_ArraySlice_l173_88_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_88_6 = {3'd0, _zz_when_ArraySlice_l173_88_7};
  assign _zz_when_ArraySlice_l173_88_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_89 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_89_1);
  assign _zz_when_ArraySlice_l165_89_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_89_1 = {2'd0, _zz_when_ArraySlice_l165_89_2};
  assign _zz_when_ArraySlice_l166_89 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_89_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_89_2);
  assign _zz_when_ArraySlice_l166_89_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_89_3);
  assign _zz_when_ArraySlice_l166_89_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_89_3 = {2'd0, _zz_when_ArraySlice_l166_89_4};
  assign _zz__zz_when_ArraySlice_l112_89 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_89 = (_zz_when_ArraySlice_l113_89_1 - _zz_when_ArraySlice_l113_89_4);
  assign _zz_when_ArraySlice_l113_89_1 = (_zz_when_ArraySlice_l113_89_2 + _zz_when_ArraySlice_l113_89_3);
  assign _zz_when_ArraySlice_l113_89_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_89_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_89_4 = {1'd0, _zz_when_ArraySlice_l112_89};
  assign _zz__zz_when_ArraySlice_l173_89 = (_zz__zz_when_ArraySlice_l173_89_1 + _zz__zz_when_ArraySlice_l173_89_2);
  assign _zz__zz_when_ArraySlice_l173_89_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_89_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_89_3 = {1'd0, _zz_when_ArraySlice_l112_89};
  assign _zz_when_ArraySlice_l118_89_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_89 = _zz_when_ArraySlice_l118_89_1[5:0];
  assign _zz_when_ArraySlice_l173_89_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_89_1 = {1'd0, _zz_when_ArraySlice_l173_89_2};
  assign _zz_when_ArraySlice_l173_89_3 = (_zz_when_ArraySlice_l173_89_4 + _zz_when_ArraySlice_l173_89_9);
  assign _zz_when_ArraySlice_l173_89_4 = (_zz_when_ArraySlice_l173_89 - _zz_when_ArraySlice_l173_89_5);
  assign _zz_when_ArraySlice_l173_89_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_89_7);
  assign _zz_when_ArraySlice_l173_89_5 = {1'd0, _zz_when_ArraySlice_l173_89_6};
  assign _zz_when_ArraySlice_l173_89_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_89_7 = {2'd0, _zz_when_ArraySlice_l173_89_8};
  assign _zz_when_ArraySlice_l173_89_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_90 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_90_1);
  assign _zz_when_ArraySlice_l165_90_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_90_1 = {1'd0, _zz_when_ArraySlice_l165_90_2};
  assign _zz_when_ArraySlice_l166_90 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_90_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_90_2);
  assign _zz_when_ArraySlice_l166_90_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_90_3);
  assign _zz_when_ArraySlice_l166_90_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_90_3 = {1'd0, _zz_when_ArraySlice_l166_90_4};
  assign _zz__zz_when_ArraySlice_l112_90 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_90 = (_zz_when_ArraySlice_l113_90_1 - _zz_when_ArraySlice_l113_90_4);
  assign _zz_when_ArraySlice_l113_90_1 = (_zz_when_ArraySlice_l113_90_2 + _zz_when_ArraySlice_l113_90_3);
  assign _zz_when_ArraySlice_l113_90_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_90_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_90_4 = {1'd0, _zz_when_ArraySlice_l112_90};
  assign _zz__zz_when_ArraySlice_l173_90 = (_zz__zz_when_ArraySlice_l173_90_1 + _zz__zz_when_ArraySlice_l173_90_2);
  assign _zz__zz_when_ArraySlice_l173_90_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_90_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_90_3 = {1'd0, _zz_when_ArraySlice_l112_90};
  assign _zz_when_ArraySlice_l118_90_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_90 = _zz_when_ArraySlice_l118_90_1[5:0];
  assign _zz_when_ArraySlice_l173_90_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_90_1 = {1'd0, _zz_when_ArraySlice_l173_90_2};
  assign _zz_when_ArraySlice_l173_90_3 = (_zz_when_ArraySlice_l173_90_4 + _zz_when_ArraySlice_l173_90_9);
  assign _zz_when_ArraySlice_l173_90_4 = (_zz_when_ArraySlice_l173_90 - _zz_when_ArraySlice_l173_90_5);
  assign _zz_when_ArraySlice_l173_90_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_90_7);
  assign _zz_when_ArraySlice_l173_90_5 = {1'd0, _zz_when_ArraySlice_l173_90_6};
  assign _zz_when_ArraySlice_l173_90_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_90_7 = {1'd0, _zz_when_ArraySlice_l173_90_8};
  assign _zz_when_ArraySlice_l173_90_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_91 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_91_1);
  assign _zz_when_ArraySlice_l165_91_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_91_1 = {1'd0, _zz_when_ArraySlice_l165_91_2};
  assign _zz_when_ArraySlice_l166_91 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_91_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_91_2);
  assign _zz_when_ArraySlice_l166_91_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_91_3);
  assign _zz_when_ArraySlice_l166_91_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_91_3 = {1'd0, _zz_when_ArraySlice_l166_91_4};
  assign _zz__zz_when_ArraySlice_l112_91 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_91 = (_zz_when_ArraySlice_l113_91_1 - _zz_when_ArraySlice_l113_91_4);
  assign _zz_when_ArraySlice_l113_91_1 = (_zz_when_ArraySlice_l113_91_2 + _zz_when_ArraySlice_l113_91_3);
  assign _zz_when_ArraySlice_l113_91_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_91_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_91_4 = {1'd0, _zz_when_ArraySlice_l112_91};
  assign _zz__zz_when_ArraySlice_l173_91 = (_zz__zz_when_ArraySlice_l173_91_1 + _zz__zz_when_ArraySlice_l173_91_2);
  assign _zz__zz_when_ArraySlice_l173_91_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_91_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_91_3 = {1'd0, _zz_when_ArraySlice_l112_91};
  assign _zz_when_ArraySlice_l118_91_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_91 = _zz_when_ArraySlice_l118_91_1[5:0];
  assign _zz_when_ArraySlice_l173_91_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_91_1 = {1'd0, _zz_when_ArraySlice_l173_91_2};
  assign _zz_when_ArraySlice_l173_91_3 = (_zz_when_ArraySlice_l173_91_4 + _zz_when_ArraySlice_l173_91_9);
  assign _zz_when_ArraySlice_l173_91_4 = (_zz_when_ArraySlice_l173_91 - _zz_when_ArraySlice_l173_91_5);
  assign _zz_when_ArraySlice_l173_91_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_91_7);
  assign _zz_when_ArraySlice_l173_91_5 = {1'd0, _zz_when_ArraySlice_l173_91_6};
  assign _zz_when_ArraySlice_l173_91_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_91_7 = {1'd0, _zz_when_ArraySlice_l173_91_8};
  assign _zz_when_ArraySlice_l173_91_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_92 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_92_1);
  assign _zz_when_ArraySlice_l165_92_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_92 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_92_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_92_2);
  assign _zz_when_ArraySlice_l166_92_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_92_3);
  assign _zz_when_ArraySlice_l166_92_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_92 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_92 = (_zz_when_ArraySlice_l113_92_1 - _zz_when_ArraySlice_l113_92_4);
  assign _zz_when_ArraySlice_l113_92_1 = (_zz_when_ArraySlice_l113_92_2 + _zz_when_ArraySlice_l113_92_3);
  assign _zz_when_ArraySlice_l113_92_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_92_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_92_4 = {1'd0, _zz_when_ArraySlice_l112_92};
  assign _zz__zz_when_ArraySlice_l173_92 = (_zz__zz_when_ArraySlice_l173_92_1 + _zz__zz_when_ArraySlice_l173_92_2);
  assign _zz__zz_when_ArraySlice_l173_92_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_92_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_92_3 = {1'd0, _zz_when_ArraySlice_l112_92};
  assign _zz_when_ArraySlice_l118_92_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_92 = _zz_when_ArraySlice_l118_92_1[5:0];
  assign _zz_when_ArraySlice_l173_92_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_92_1 = {1'd0, _zz_when_ArraySlice_l173_92_2};
  assign _zz_when_ArraySlice_l173_92_3 = (_zz_when_ArraySlice_l173_92_4 + _zz_when_ArraySlice_l173_92_8);
  assign _zz_when_ArraySlice_l173_92_4 = (_zz_when_ArraySlice_l173_92 - _zz_when_ArraySlice_l173_92_5);
  assign _zz_when_ArraySlice_l173_92_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_92_7);
  assign _zz_when_ArraySlice_l173_92_5 = {1'd0, _zz_when_ArraySlice_l173_92_6};
  assign _zz_when_ArraySlice_l173_92_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_92_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_93 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_93_1);
  assign _zz_when_ArraySlice_l165_93_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_93_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_93 = {1'd0, _zz_when_ArraySlice_l166_93_1};
  assign _zz_when_ArraySlice_l166_93_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_93_3);
  assign _zz_when_ArraySlice_l166_93_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_93_4);
  assign _zz_when_ArraySlice_l166_93_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_93 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_93 = (_zz_when_ArraySlice_l113_93_1 - _zz_when_ArraySlice_l113_93_4);
  assign _zz_when_ArraySlice_l113_93_1 = (_zz_when_ArraySlice_l113_93_2 + _zz_when_ArraySlice_l113_93_3);
  assign _zz_when_ArraySlice_l113_93_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_93_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_93_4 = {1'd0, _zz_when_ArraySlice_l112_93};
  assign _zz__zz_when_ArraySlice_l173_93 = (_zz__zz_when_ArraySlice_l173_93_1 + _zz__zz_when_ArraySlice_l173_93_2);
  assign _zz__zz_when_ArraySlice_l173_93_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_93_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_93_3 = {1'd0, _zz_when_ArraySlice_l112_93};
  assign _zz_when_ArraySlice_l118_93_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_93 = _zz_when_ArraySlice_l118_93_1[5:0];
  assign _zz_when_ArraySlice_l173_93_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_93_1 = {2'd0, _zz_when_ArraySlice_l173_93_2};
  assign _zz_when_ArraySlice_l173_93_3 = (_zz_when_ArraySlice_l173_93_4 + _zz_when_ArraySlice_l173_93_8);
  assign _zz_when_ArraySlice_l173_93_4 = (_zz_when_ArraySlice_l173_93 - _zz_when_ArraySlice_l173_93_5);
  assign _zz_when_ArraySlice_l173_93_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_93_7);
  assign _zz_when_ArraySlice_l173_93_5 = {1'd0, _zz_when_ArraySlice_l173_93_6};
  assign _zz_when_ArraySlice_l173_93_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_93_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_94 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_94_1);
  assign _zz_when_ArraySlice_l165_94_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_94_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_94 = {1'd0, _zz_when_ArraySlice_l166_94_1};
  assign _zz_when_ArraySlice_l166_94_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_94_3);
  assign _zz_when_ArraySlice_l166_94_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_94_4);
  assign _zz_when_ArraySlice_l166_94_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_94 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_94 = (_zz_when_ArraySlice_l113_94_1 - _zz_when_ArraySlice_l113_94_4);
  assign _zz_when_ArraySlice_l113_94_1 = (_zz_when_ArraySlice_l113_94_2 + _zz_when_ArraySlice_l113_94_3);
  assign _zz_when_ArraySlice_l113_94_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_94_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_94_4 = {1'd0, _zz_when_ArraySlice_l112_94};
  assign _zz__zz_when_ArraySlice_l173_94 = (_zz__zz_when_ArraySlice_l173_94_1 + _zz__zz_when_ArraySlice_l173_94_2);
  assign _zz__zz_when_ArraySlice_l173_94_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_94_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_94_3 = {1'd0, _zz_when_ArraySlice_l112_94};
  assign _zz_when_ArraySlice_l118_94_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_94 = _zz_when_ArraySlice_l118_94_1[5:0];
  assign _zz_when_ArraySlice_l173_94_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_94_1 = {2'd0, _zz_when_ArraySlice_l173_94_2};
  assign _zz_when_ArraySlice_l173_94_3 = (_zz_when_ArraySlice_l173_94_4 + _zz_when_ArraySlice_l173_94_8);
  assign _zz_when_ArraySlice_l173_94_4 = (_zz_when_ArraySlice_l173_94 - _zz_when_ArraySlice_l173_94_5);
  assign _zz_when_ArraySlice_l173_94_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_94_7);
  assign _zz_when_ArraySlice_l173_94_5 = {1'd0, _zz_when_ArraySlice_l173_94_6};
  assign _zz_when_ArraySlice_l173_94_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_94_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_95 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_95_1);
  assign _zz_when_ArraySlice_l165_95_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_95_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_95 = {2'd0, _zz_when_ArraySlice_l166_95_1};
  assign _zz_when_ArraySlice_l166_95_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_95_3);
  assign _zz_when_ArraySlice_l166_95_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_95_4);
  assign _zz_when_ArraySlice_l166_95_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_95 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_95 = (_zz_when_ArraySlice_l113_95_1 - _zz_when_ArraySlice_l113_95_4);
  assign _zz_when_ArraySlice_l113_95_1 = (_zz_when_ArraySlice_l113_95_2 + _zz_when_ArraySlice_l113_95_3);
  assign _zz_when_ArraySlice_l113_95_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_95_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_95_4 = {1'd0, _zz_when_ArraySlice_l112_95};
  assign _zz__zz_when_ArraySlice_l173_95 = (_zz__zz_when_ArraySlice_l173_95_1 + _zz__zz_when_ArraySlice_l173_95_2);
  assign _zz__zz_when_ArraySlice_l173_95_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_95_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_95_3 = {1'd0, _zz_when_ArraySlice_l112_95};
  assign _zz_when_ArraySlice_l118_95_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_95 = _zz_when_ArraySlice_l118_95_1[5:0];
  assign _zz_when_ArraySlice_l173_95_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_95_1 = {3'd0, _zz_when_ArraySlice_l173_95_2};
  assign _zz_when_ArraySlice_l173_95_3 = (_zz_when_ArraySlice_l173_95_4 + _zz_when_ArraySlice_l173_95_8);
  assign _zz_when_ArraySlice_l173_95_4 = (_zz_when_ArraySlice_l173_95 - _zz_when_ArraySlice_l173_95_5);
  assign _zz_when_ArraySlice_l173_95_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_95_7);
  assign _zz_when_ArraySlice_l173_95_5 = {1'd0, _zz_when_ArraySlice_l173_95_6};
  assign _zz_when_ArraySlice_l173_95_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_95_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l421_3_1 = (_zz_when_ArraySlice_l421_3_2 + _zz_when_ArraySlice_l421_3_7);
  assign _zz_when_ArraySlice_l421_3_2 = (_zz_when_ArraySlice_l421_3_3 + _zz_when_ArraySlice_l421_3_5);
  assign _zz_when_ArraySlice_l421_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l421_3_4);
  assign _zz_when_ArraySlice_l421_3_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l421_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l421_3_5 = {5'd0, _zz_when_ArraySlice_l421_3_6};
  assign _zz_when_ArraySlice_l421_3_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l421_3_7 = {1'd0, _zz_when_ArraySlice_l421_3_8};
  assign _zz_selectReadFifo_3_25 = 1'b1;
  assign _zz_selectReadFifo_3_24 = {5'd0, _zz_selectReadFifo_3_25};
  assign _zz_when_ArraySlice_l425_3_1 = (_zz_when_ArraySlice_l425_3_2 % aReg);
  assign _zz_when_ArraySlice_l425_3_2 = (handshakeTimes_3_value + _zz_when_ArraySlice_l425_3_3);
  assign _zz_when_ArraySlice_l425_3_4 = 1'b1;
  assign _zz_when_ArraySlice_l425_3_3 = {12'd0, _zz_when_ArraySlice_l425_3_4};
  assign _zz_when_ArraySlice_l436_3_2 = (_zz_when_ArraySlice_l436_3_3 - _zz_when_ArraySlice_l436_3_4);
  assign _zz_when_ArraySlice_l436_3_1 = {7'd0, _zz_when_ArraySlice_l436_3_2};
  assign _zz_when_ArraySlice_l436_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l436_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l436_3_4 = {5'd0, _zz_when_ArraySlice_l436_3_5};
  assign _zz__zz_when_ArraySlice_l94_11 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_11 = (_zz_when_ArraySlice_l95_11_1 - _zz_when_ArraySlice_l95_11_4);
  assign _zz_when_ArraySlice_l95_11_1 = (_zz_when_ArraySlice_l95_11_2 + _zz_when_ArraySlice_l95_11_3);
  assign _zz_when_ArraySlice_l95_11_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_11_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_11_4 = {1'd0, _zz_when_ArraySlice_l94_11};
  assign _zz__zz_when_ArraySlice_l437_3_1 = (_zz__zz_when_ArraySlice_l437_3_2 + _zz__zz_when_ArraySlice_l437_3_3);
  assign _zz__zz_when_ArraySlice_l437_3_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l437_3_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l437_3_4 = {1'd0, _zz_when_ArraySlice_l94_11};
  assign _zz_when_ArraySlice_l99_11_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_11 = _zz_when_ArraySlice_l99_11_1[5:0];
  assign _zz_when_ArraySlice_l437_3_1 = (outSliceNumb_3_value + _zz_when_ArraySlice_l437_3_2);
  assign _zz_when_ArraySlice_l437_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l437_3_2 = {6'd0, _zz_when_ArraySlice_l437_3_3};
  assign _zz_when_ArraySlice_l437_3_4 = (_zz_when_ArraySlice_l437_3 / aReg);
  assign _zz_selectReadFifo_3_26 = (selectReadFifo_3 - _zz_selectReadFifo_3_27);
  assign _zz_selectReadFifo_3_27 = {3'd0, bReg};
  assign _zz_selectReadFifo_3_29 = 1'b1;
  assign _zz_selectReadFifo_3_28 = {5'd0, _zz_selectReadFifo_3_29};
  assign _zz_when_ArraySlice_l165_96 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_96_1);
  assign _zz_when_ArraySlice_l165_96_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_96_1 = {3'd0, _zz_when_ArraySlice_l165_96_2};
  assign _zz_when_ArraySlice_l166_96 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_96_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_96_3);
  assign _zz_when_ArraySlice_l166_96_1 = {1'd0, _zz_when_ArraySlice_l166_96_2};
  assign _zz_when_ArraySlice_l166_96_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_96_4);
  assign _zz_when_ArraySlice_l166_96_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_96_4 = {3'd0, _zz_when_ArraySlice_l166_96_5};
  assign _zz__zz_when_ArraySlice_l112_96 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_96 = (_zz_when_ArraySlice_l113_96_1 - _zz_when_ArraySlice_l113_96_4);
  assign _zz_when_ArraySlice_l113_96_1 = (_zz_when_ArraySlice_l113_96_2 + _zz_when_ArraySlice_l113_96_3);
  assign _zz_when_ArraySlice_l113_96_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_96_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_96_4 = {1'd0, _zz_when_ArraySlice_l112_96};
  assign _zz__zz_when_ArraySlice_l173_96 = (_zz__zz_when_ArraySlice_l173_96_1 + _zz__zz_when_ArraySlice_l173_96_2);
  assign _zz__zz_when_ArraySlice_l173_96_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_96_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_96_3 = {1'd0, _zz_when_ArraySlice_l112_96};
  assign _zz_when_ArraySlice_l118_96_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_96 = _zz_when_ArraySlice_l118_96_1[5:0];
  assign _zz_when_ArraySlice_l173_96_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_96_2 = (_zz_when_ArraySlice_l173_96_3 + _zz_when_ArraySlice_l173_96_8);
  assign _zz_when_ArraySlice_l173_96_3 = (_zz_when_ArraySlice_l173_96 - _zz_when_ArraySlice_l173_96_4);
  assign _zz_when_ArraySlice_l173_96_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_96_6);
  assign _zz_when_ArraySlice_l173_96_4 = {1'd0, _zz_when_ArraySlice_l173_96_5};
  assign _zz_when_ArraySlice_l173_96_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_96_6 = {3'd0, _zz_when_ArraySlice_l173_96_7};
  assign _zz_when_ArraySlice_l173_96_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_97 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_97_1);
  assign _zz_when_ArraySlice_l165_97_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_97_1 = {2'd0, _zz_when_ArraySlice_l165_97_2};
  assign _zz_when_ArraySlice_l166_97 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_97_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_97_2);
  assign _zz_when_ArraySlice_l166_97_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_97_3);
  assign _zz_when_ArraySlice_l166_97_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_97_3 = {2'd0, _zz_when_ArraySlice_l166_97_4};
  assign _zz__zz_when_ArraySlice_l112_97 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_97 = (_zz_when_ArraySlice_l113_97_1 - _zz_when_ArraySlice_l113_97_4);
  assign _zz_when_ArraySlice_l113_97_1 = (_zz_when_ArraySlice_l113_97_2 + _zz_when_ArraySlice_l113_97_3);
  assign _zz_when_ArraySlice_l113_97_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_97_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_97_4 = {1'd0, _zz_when_ArraySlice_l112_97};
  assign _zz__zz_when_ArraySlice_l173_97 = (_zz__zz_when_ArraySlice_l173_97_1 + _zz__zz_when_ArraySlice_l173_97_2);
  assign _zz__zz_when_ArraySlice_l173_97_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_97_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_97_3 = {1'd0, _zz_when_ArraySlice_l112_97};
  assign _zz_when_ArraySlice_l118_97_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_97 = _zz_when_ArraySlice_l118_97_1[5:0];
  assign _zz_when_ArraySlice_l173_97_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_97_1 = {1'd0, _zz_when_ArraySlice_l173_97_2};
  assign _zz_when_ArraySlice_l173_97_3 = (_zz_when_ArraySlice_l173_97_4 + _zz_when_ArraySlice_l173_97_9);
  assign _zz_when_ArraySlice_l173_97_4 = (_zz_when_ArraySlice_l173_97 - _zz_when_ArraySlice_l173_97_5);
  assign _zz_when_ArraySlice_l173_97_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_97_7);
  assign _zz_when_ArraySlice_l173_97_5 = {1'd0, _zz_when_ArraySlice_l173_97_6};
  assign _zz_when_ArraySlice_l173_97_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_97_7 = {2'd0, _zz_when_ArraySlice_l173_97_8};
  assign _zz_when_ArraySlice_l173_97_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_98 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_98_1);
  assign _zz_when_ArraySlice_l165_98_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_98_1 = {1'd0, _zz_when_ArraySlice_l165_98_2};
  assign _zz_when_ArraySlice_l166_98 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_98_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_98_2);
  assign _zz_when_ArraySlice_l166_98_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_98_3);
  assign _zz_when_ArraySlice_l166_98_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_98_3 = {1'd0, _zz_when_ArraySlice_l166_98_4};
  assign _zz__zz_when_ArraySlice_l112_98 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_98 = (_zz_when_ArraySlice_l113_98_1 - _zz_when_ArraySlice_l113_98_4);
  assign _zz_when_ArraySlice_l113_98_1 = (_zz_when_ArraySlice_l113_98_2 + _zz_when_ArraySlice_l113_98_3);
  assign _zz_when_ArraySlice_l113_98_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_98_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_98_4 = {1'd0, _zz_when_ArraySlice_l112_98};
  assign _zz__zz_when_ArraySlice_l173_98 = (_zz__zz_when_ArraySlice_l173_98_1 + _zz__zz_when_ArraySlice_l173_98_2);
  assign _zz__zz_when_ArraySlice_l173_98_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_98_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_98_3 = {1'd0, _zz_when_ArraySlice_l112_98};
  assign _zz_when_ArraySlice_l118_98_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_98 = _zz_when_ArraySlice_l118_98_1[5:0];
  assign _zz_when_ArraySlice_l173_98_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_98_1 = {1'd0, _zz_when_ArraySlice_l173_98_2};
  assign _zz_when_ArraySlice_l173_98_3 = (_zz_when_ArraySlice_l173_98_4 + _zz_when_ArraySlice_l173_98_9);
  assign _zz_when_ArraySlice_l173_98_4 = (_zz_when_ArraySlice_l173_98 - _zz_when_ArraySlice_l173_98_5);
  assign _zz_when_ArraySlice_l173_98_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_98_7);
  assign _zz_when_ArraySlice_l173_98_5 = {1'd0, _zz_when_ArraySlice_l173_98_6};
  assign _zz_when_ArraySlice_l173_98_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_98_7 = {1'd0, _zz_when_ArraySlice_l173_98_8};
  assign _zz_when_ArraySlice_l173_98_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_99 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_99_1);
  assign _zz_when_ArraySlice_l165_99_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_99_1 = {1'd0, _zz_when_ArraySlice_l165_99_2};
  assign _zz_when_ArraySlice_l166_99 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_99_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_99_2);
  assign _zz_when_ArraySlice_l166_99_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_99_3);
  assign _zz_when_ArraySlice_l166_99_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_99_3 = {1'd0, _zz_when_ArraySlice_l166_99_4};
  assign _zz__zz_when_ArraySlice_l112_99 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_99 = (_zz_when_ArraySlice_l113_99_1 - _zz_when_ArraySlice_l113_99_4);
  assign _zz_when_ArraySlice_l113_99_1 = (_zz_when_ArraySlice_l113_99_2 + _zz_when_ArraySlice_l113_99_3);
  assign _zz_when_ArraySlice_l113_99_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_99_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_99_4 = {1'd0, _zz_when_ArraySlice_l112_99};
  assign _zz__zz_when_ArraySlice_l173_99 = (_zz__zz_when_ArraySlice_l173_99_1 + _zz__zz_when_ArraySlice_l173_99_2);
  assign _zz__zz_when_ArraySlice_l173_99_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_99_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_99_3 = {1'd0, _zz_when_ArraySlice_l112_99};
  assign _zz_when_ArraySlice_l118_99_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_99 = _zz_when_ArraySlice_l118_99_1[5:0];
  assign _zz_when_ArraySlice_l173_99_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_99_1 = {1'd0, _zz_when_ArraySlice_l173_99_2};
  assign _zz_when_ArraySlice_l173_99_3 = (_zz_when_ArraySlice_l173_99_4 + _zz_when_ArraySlice_l173_99_9);
  assign _zz_when_ArraySlice_l173_99_4 = (_zz_when_ArraySlice_l173_99 - _zz_when_ArraySlice_l173_99_5);
  assign _zz_when_ArraySlice_l173_99_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_99_7);
  assign _zz_when_ArraySlice_l173_99_5 = {1'd0, _zz_when_ArraySlice_l173_99_6};
  assign _zz_when_ArraySlice_l173_99_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_99_7 = {1'd0, _zz_when_ArraySlice_l173_99_8};
  assign _zz_when_ArraySlice_l173_99_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_100 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_100_1);
  assign _zz_when_ArraySlice_l165_100_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_100 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_100_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_100_2);
  assign _zz_when_ArraySlice_l166_100_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_100_3);
  assign _zz_when_ArraySlice_l166_100_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_100 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_100 = (_zz_when_ArraySlice_l113_100_1 - _zz_when_ArraySlice_l113_100_4);
  assign _zz_when_ArraySlice_l113_100_1 = (_zz_when_ArraySlice_l113_100_2 + _zz_when_ArraySlice_l113_100_3);
  assign _zz_when_ArraySlice_l113_100_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_100_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_100_4 = {1'd0, _zz_when_ArraySlice_l112_100};
  assign _zz__zz_when_ArraySlice_l173_100 = (_zz__zz_when_ArraySlice_l173_100_1 + _zz__zz_when_ArraySlice_l173_100_2);
  assign _zz__zz_when_ArraySlice_l173_100_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_100_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_100_3 = {1'd0, _zz_when_ArraySlice_l112_100};
  assign _zz_when_ArraySlice_l118_100_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_100 = _zz_when_ArraySlice_l118_100_1[5:0];
  assign _zz_when_ArraySlice_l173_100_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_100_1 = {1'd0, _zz_when_ArraySlice_l173_100_2};
  assign _zz_when_ArraySlice_l173_100_3 = (_zz_when_ArraySlice_l173_100_4 + _zz_when_ArraySlice_l173_100_8);
  assign _zz_when_ArraySlice_l173_100_4 = (_zz_when_ArraySlice_l173_100 - _zz_when_ArraySlice_l173_100_5);
  assign _zz_when_ArraySlice_l173_100_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_100_7);
  assign _zz_when_ArraySlice_l173_100_5 = {1'd0, _zz_when_ArraySlice_l173_100_6};
  assign _zz_when_ArraySlice_l173_100_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_100_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_101 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_101_1);
  assign _zz_when_ArraySlice_l165_101_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_101_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_101 = {1'd0, _zz_when_ArraySlice_l166_101_1};
  assign _zz_when_ArraySlice_l166_101_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_101_3);
  assign _zz_when_ArraySlice_l166_101_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_101_4);
  assign _zz_when_ArraySlice_l166_101_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_101 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_101 = (_zz_when_ArraySlice_l113_101_1 - _zz_when_ArraySlice_l113_101_4);
  assign _zz_when_ArraySlice_l113_101_1 = (_zz_when_ArraySlice_l113_101_2 + _zz_when_ArraySlice_l113_101_3);
  assign _zz_when_ArraySlice_l113_101_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_101_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_101_4 = {1'd0, _zz_when_ArraySlice_l112_101};
  assign _zz__zz_when_ArraySlice_l173_101 = (_zz__zz_when_ArraySlice_l173_101_1 + _zz__zz_when_ArraySlice_l173_101_2);
  assign _zz__zz_when_ArraySlice_l173_101_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_101_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_101_3 = {1'd0, _zz_when_ArraySlice_l112_101};
  assign _zz_when_ArraySlice_l118_101_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_101 = _zz_when_ArraySlice_l118_101_1[5:0];
  assign _zz_when_ArraySlice_l173_101_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_101_1 = {2'd0, _zz_when_ArraySlice_l173_101_2};
  assign _zz_when_ArraySlice_l173_101_3 = (_zz_when_ArraySlice_l173_101_4 + _zz_when_ArraySlice_l173_101_8);
  assign _zz_when_ArraySlice_l173_101_4 = (_zz_when_ArraySlice_l173_101 - _zz_when_ArraySlice_l173_101_5);
  assign _zz_when_ArraySlice_l173_101_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_101_7);
  assign _zz_when_ArraySlice_l173_101_5 = {1'd0, _zz_when_ArraySlice_l173_101_6};
  assign _zz_when_ArraySlice_l173_101_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_101_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_102 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_102_1);
  assign _zz_when_ArraySlice_l165_102_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_102_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_102 = {1'd0, _zz_when_ArraySlice_l166_102_1};
  assign _zz_when_ArraySlice_l166_102_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_102_3);
  assign _zz_when_ArraySlice_l166_102_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_102_4);
  assign _zz_when_ArraySlice_l166_102_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_102 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_102 = (_zz_when_ArraySlice_l113_102_1 - _zz_when_ArraySlice_l113_102_4);
  assign _zz_when_ArraySlice_l113_102_1 = (_zz_when_ArraySlice_l113_102_2 + _zz_when_ArraySlice_l113_102_3);
  assign _zz_when_ArraySlice_l113_102_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_102_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_102_4 = {1'd0, _zz_when_ArraySlice_l112_102};
  assign _zz__zz_when_ArraySlice_l173_102 = (_zz__zz_when_ArraySlice_l173_102_1 + _zz__zz_when_ArraySlice_l173_102_2);
  assign _zz__zz_when_ArraySlice_l173_102_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_102_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_102_3 = {1'd0, _zz_when_ArraySlice_l112_102};
  assign _zz_when_ArraySlice_l118_102_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_102 = _zz_when_ArraySlice_l118_102_1[5:0];
  assign _zz_when_ArraySlice_l173_102_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_102_1 = {2'd0, _zz_when_ArraySlice_l173_102_2};
  assign _zz_when_ArraySlice_l173_102_3 = (_zz_when_ArraySlice_l173_102_4 + _zz_when_ArraySlice_l173_102_8);
  assign _zz_when_ArraySlice_l173_102_4 = (_zz_when_ArraySlice_l173_102 - _zz_when_ArraySlice_l173_102_5);
  assign _zz_when_ArraySlice_l173_102_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_102_7);
  assign _zz_when_ArraySlice_l173_102_5 = {1'd0, _zz_when_ArraySlice_l173_102_6};
  assign _zz_when_ArraySlice_l173_102_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_102_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_103 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_103_1);
  assign _zz_when_ArraySlice_l165_103_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_103_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_103 = {2'd0, _zz_when_ArraySlice_l166_103_1};
  assign _zz_when_ArraySlice_l166_103_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_103_3);
  assign _zz_when_ArraySlice_l166_103_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_103_4);
  assign _zz_when_ArraySlice_l166_103_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_103 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_103 = (_zz_when_ArraySlice_l113_103_1 - _zz_when_ArraySlice_l113_103_4);
  assign _zz_when_ArraySlice_l113_103_1 = (_zz_when_ArraySlice_l113_103_2 + _zz_when_ArraySlice_l113_103_3);
  assign _zz_when_ArraySlice_l113_103_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_103_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_103_4 = {1'd0, _zz_when_ArraySlice_l112_103};
  assign _zz__zz_when_ArraySlice_l173_103 = (_zz__zz_when_ArraySlice_l173_103_1 + _zz__zz_when_ArraySlice_l173_103_2);
  assign _zz__zz_when_ArraySlice_l173_103_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_103_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_103_3 = {1'd0, _zz_when_ArraySlice_l112_103};
  assign _zz_when_ArraySlice_l118_103_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_103 = _zz_when_ArraySlice_l118_103_1[5:0];
  assign _zz_when_ArraySlice_l173_103_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_103_1 = {3'd0, _zz_when_ArraySlice_l173_103_2};
  assign _zz_when_ArraySlice_l173_103_3 = (_zz_when_ArraySlice_l173_103_4 + _zz_when_ArraySlice_l173_103_8);
  assign _zz_when_ArraySlice_l173_103_4 = (_zz_when_ArraySlice_l173_103 - _zz_when_ArraySlice_l173_103_5);
  assign _zz_when_ArraySlice_l173_103_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_103_7);
  assign _zz_when_ArraySlice_l173_103_5 = {1'd0, _zz_when_ArraySlice_l173_103_6};
  assign _zz_when_ArraySlice_l173_103_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_103_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_3_31 = 1'b1;
  assign _zz_selectReadFifo_3_30 = {5'd0, _zz_selectReadFifo_3_31};
  assign _zz_when_ArraySlice_l448_3_1 = (_zz_when_ArraySlice_l448_3_2 % aReg);
  assign _zz_when_ArraySlice_l448_3_2 = (handshakeTimes_3_value + _zz_when_ArraySlice_l448_3_3);
  assign _zz_when_ArraySlice_l448_3_4 = 1'b1;
  assign _zz_when_ArraySlice_l448_3_3 = {12'd0, _zz_when_ArraySlice_l448_3_4};
  assign _zz_when_ArraySlice_l434_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l434_3_1);
  assign _zz_when_ArraySlice_l434_3_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l434_3_1 = {1'd0, _zz_when_ArraySlice_l434_3_2};
  assign _zz_when_ArraySlice_l455_3_2 = (_zz_when_ArraySlice_l455_3_3 - _zz_when_ArraySlice_l455_3_4);
  assign _zz_when_ArraySlice_l455_3_1 = {7'd0, _zz_when_ArraySlice_l455_3_2};
  assign _zz_when_ArraySlice_l455_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l455_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l455_3_4 = {5'd0, _zz_when_ArraySlice_l455_3_5};
  assign _zz_when_ArraySlice_l373_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l373_4_1);
  assign _zz_when_ArraySlice_l373_4_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l374_4_1 = (selectReadFifo_4 + _zz_when_ArraySlice_l374_4_2);
  assign _zz_when_ArraySlice_l374_4_2 = (bReg * 3'b100);
  assign _zz__zz_outputStreamArrayData_4_valid = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l380_4_2 = 1'b1;
  assign _zz_when_ArraySlice_l380_4_1 = {6'd0, _zz_when_ArraySlice_l380_4_2};
  assign _zz_when_ArraySlice_l380_4_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l380_4_5);
  assign _zz_when_ArraySlice_l380_4_5 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l381_4_2 = (_zz_when_ArraySlice_l381_4_3 - _zz_when_ArraySlice_l381_4_4);
  assign _zz_when_ArraySlice_l381_4_1 = {7'd0, _zz_when_ArraySlice_l381_4_2};
  assign _zz_when_ArraySlice_l381_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l381_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l381_4_4 = {5'd0, _zz_when_ArraySlice_l381_4_5};
  assign _zz_selectReadFifo_4 = (selectReadFifo_4 - _zz_selectReadFifo_4_1);
  assign _zz_selectReadFifo_4_1 = {3'd0, bReg};
  assign _zz_selectReadFifo_4_3 = 1'b1;
  assign _zz_selectReadFifo_4_2 = {5'd0, _zz_selectReadFifo_4_3};
  assign _zz_selectReadFifo_4_5 = 1'b1;
  assign _zz_selectReadFifo_4_4 = {5'd0, _zz_selectReadFifo_4_5};
  assign _zz_when_ArraySlice_l384_4 = (_zz_when_ArraySlice_l384_4_1 % aReg);
  assign _zz_when_ArraySlice_l384_4_1 = (handshakeTimes_4_value + _zz_when_ArraySlice_l384_4_2);
  assign _zz_when_ArraySlice_l384_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l384_4_2 = {12'd0, _zz_when_ArraySlice_l384_4_3};
  assign _zz_when_ArraySlice_l389_4_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l389_4_3);
  assign _zz_when_ArraySlice_l389_4_3 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l389_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l389_4_4 = {6'd0, _zz_when_ArraySlice_l389_4_5};
  assign _zz_when_ArraySlice_l390_4_2 = (_zz_when_ArraySlice_l390_4_3 - _zz_when_ArraySlice_l390_4_4);
  assign _zz_when_ArraySlice_l390_4_1 = {7'd0, _zz_when_ArraySlice_l390_4_2};
  assign _zz_when_ArraySlice_l390_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l390_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l390_4_4 = {5'd0, _zz_when_ArraySlice_l390_4_5};
  assign _zz__zz_when_ArraySlice_l94_12 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_12 = (_zz_when_ArraySlice_l95_12_1 - _zz_when_ArraySlice_l95_12_4);
  assign _zz_when_ArraySlice_l95_12_1 = (_zz_when_ArraySlice_l95_12_2 + _zz_when_ArraySlice_l95_12_3);
  assign _zz_when_ArraySlice_l95_12_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_12_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_12_4 = {1'd0, _zz_when_ArraySlice_l94_12};
  assign _zz__zz_when_ArraySlice_l392_4 = (_zz__zz_when_ArraySlice_l392_4_1 + _zz__zz_when_ArraySlice_l392_4_2);
  assign _zz__zz_when_ArraySlice_l392_4_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l392_4_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l392_4_3 = {1'd0, _zz_when_ArraySlice_l94_12};
  assign _zz_when_ArraySlice_l99_12_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_12 = _zz_when_ArraySlice_l99_12_1[5:0];
  assign _zz_when_ArraySlice_l392_4_1 = (outSliceNumb_4_value + _zz_when_ArraySlice_l392_4_2);
  assign _zz_when_ArraySlice_l392_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l392_4_2 = {6'd0, _zz_when_ArraySlice_l392_4_3};
  assign _zz_when_ArraySlice_l392_4_4 = (_zz_when_ArraySlice_l392_4 / aReg);
  assign _zz_selectReadFifo_4_6 = (selectReadFifo_4 - _zz_selectReadFifo_4_7);
  assign _zz_selectReadFifo_4_7 = {3'd0, bReg};
  assign _zz_selectReadFifo_4_9 = 1'b1;
  assign _zz_selectReadFifo_4_8 = {5'd0, _zz_selectReadFifo_4_9};
  assign _zz_selectReadFifo_4_10 = (selectReadFifo_4 + _zz_selectReadFifo_4_11);
  assign _zz_selectReadFifo_4_11 = (3'b111 * bReg);
  assign _zz_selectReadFifo_4_13 = 1'b1;
  assign _zz_selectReadFifo_4_12 = {5'd0, _zz_selectReadFifo_4_13};
  assign _zz_when_ArraySlice_l165_104 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_104_1);
  assign _zz_when_ArraySlice_l165_104_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_104_1 = {3'd0, _zz_when_ArraySlice_l165_104_2};
  assign _zz_when_ArraySlice_l166_104 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_104_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_104_3);
  assign _zz_when_ArraySlice_l166_104_1 = {1'd0, _zz_when_ArraySlice_l166_104_2};
  assign _zz_when_ArraySlice_l166_104_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_104_4);
  assign _zz_when_ArraySlice_l166_104_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_104_4 = {3'd0, _zz_when_ArraySlice_l166_104_5};
  assign _zz__zz_when_ArraySlice_l112_104 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_104 = (_zz_when_ArraySlice_l113_104_1 - _zz_when_ArraySlice_l113_104_4);
  assign _zz_when_ArraySlice_l113_104_1 = (_zz_when_ArraySlice_l113_104_2 + _zz_when_ArraySlice_l113_104_3);
  assign _zz_when_ArraySlice_l113_104_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_104_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_104_4 = {1'd0, _zz_when_ArraySlice_l112_104};
  assign _zz__zz_when_ArraySlice_l173_104 = (_zz__zz_when_ArraySlice_l173_104_1 + _zz__zz_when_ArraySlice_l173_104_2);
  assign _zz__zz_when_ArraySlice_l173_104_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_104_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_104_3 = {1'd0, _zz_when_ArraySlice_l112_104};
  assign _zz_when_ArraySlice_l118_104_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_104 = _zz_when_ArraySlice_l118_104_1[5:0];
  assign _zz_when_ArraySlice_l173_104_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_104_2 = (_zz_when_ArraySlice_l173_104_3 + _zz_when_ArraySlice_l173_104_8);
  assign _zz_when_ArraySlice_l173_104_3 = (_zz_when_ArraySlice_l173_104 - _zz_when_ArraySlice_l173_104_4);
  assign _zz_when_ArraySlice_l173_104_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_104_6);
  assign _zz_when_ArraySlice_l173_104_4 = {1'd0, _zz_when_ArraySlice_l173_104_5};
  assign _zz_when_ArraySlice_l173_104_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_104_6 = {3'd0, _zz_when_ArraySlice_l173_104_7};
  assign _zz_when_ArraySlice_l173_104_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_105 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_105_1);
  assign _zz_when_ArraySlice_l165_105_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_105_1 = {2'd0, _zz_when_ArraySlice_l165_105_2};
  assign _zz_when_ArraySlice_l166_105 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_105_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_105_2);
  assign _zz_when_ArraySlice_l166_105_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_105_3);
  assign _zz_when_ArraySlice_l166_105_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_105_3 = {2'd0, _zz_when_ArraySlice_l166_105_4};
  assign _zz__zz_when_ArraySlice_l112_105 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_105 = (_zz_when_ArraySlice_l113_105_1 - _zz_when_ArraySlice_l113_105_4);
  assign _zz_when_ArraySlice_l113_105_1 = (_zz_when_ArraySlice_l113_105_2 + _zz_when_ArraySlice_l113_105_3);
  assign _zz_when_ArraySlice_l113_105_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_105_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_105_4 = {1'd0, _zz_when_ArraySlice_l112_105};
  assign _zz__zz_when_ArraySlice_l173_105 = (_zz__zz_when_ArraySlice_l173_105_1 + _zz__zz_when_ArraySlice_l173_105_2);
  assign _zz__zz_when_ArraySlice_l173_105_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_105_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_105_3 = {1'd0, _zz_when_ArraySlice_l112_105};
  assign _zz_when_ArraySlice_l118_105_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_105 = _zz_when_ArraySlice_l118_105_1[5:0];
  assign _zz_when_ArraySlice_l173_105_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_105_1 = {1'd0, _zz_when_ArraySlice_l173_105_2};
  assign _zz_when_ArraySlice_l173_105_3 = (_zz_when_ArraySlice_l173_105_4 + _zz_when_ArraySlice_l173_105_9);
  assign _zz_when_ArraySlice_l173_105_4 = (_zz_when_ArraySlice_l173_105 - _zz_when_ArraySlice_l173_105_5);
  assign _zz_when_ArraySlice_l173_105_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_105_7);
  assign _zz_when_ArraySlice_l173_105_5 = {1'd0, _zz_when_ArraySlice_l173_105_6};
  assign _zz_when_ArraySlice_l173_105_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_105_7 = {2'd0, _zz_when_ArraySlice_l173_105_8};
  assign _zz_when_ArraySlice_l173_105_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_106 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_106_1);
  assign _zz_when_ArraySlice_l165_106_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_106_1 = {1'd0, _zz_when_ArraySlice_l165_106_2};
  assign _zz_when_ArraySlice_l166_106 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_106_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_106_2);
  assign _zz_when_ArraySlice_l166_106_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_106_3);
  assign _zz_when_ArraySlice_l166_106_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_106_3 = {1'd0, _zz_when_ArraySlice_l166_106_4};
  assign _zz__zz_when_ArraySlice_l112_106 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_106 = (_zz_when_ArraySlice_l113_106_1 - _zz_when_ArraySlice_l113_106_4);
  assign _zz_when_ArraySlice_l113_106_1 = (_zz_when_ArraySlice_l113_106_2 + _zz_when_ArraySlice_l113_106_3);
  assign _zz_when_ArraySlice_l113_106_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_106_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_106_4 = {1'd0, _zz_when_ArraySlice_l112_106};
  assign _zz__zz_when_ArraySlice_l173_106 = (_zz__zz_when_ArraySlice_l173_106_1 + _zz__zz_when_ArraySlice_l173_106_2);
  assign _zz__zz_when_ArraySlice_l173_106_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_106_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_106_3 = {1'd0, _zz_when_ArraySlice_l112_106};
  assign _zz_when_ArraySlice_l118_106_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_106 = _zz_when_ArraySlice_l118_106_1[5:0];
  assign _zz_when_ArraySlice_l173_106_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_106_1 = {1'd0, _zz_when_ArraySlice_l173_106_2};
  assign _zz_when_ArraySlice_l173_106_3 = (_zz_when_ArraySlice_l173_106_4 + _zz_when_ArraySlice_l173_106_9);
  assign _zz_when_ArraySlice_l173_106_4 = (_zz_when_ArraySlice_l173_106 - _zz_when_ArraySlice_l173_106_5);
  assign _zz_when_ArraySlice_l173_106_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_106_7);
  assign _zz_when_ArraySlice_l173_106_5 = {1'd0, _zz_when_ArraySlice_l173_106_6};
  assign _zz_when_ArraySlice_l173_106_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_106_7 = {1'd0, _zz_when_ArraySlice_l173_106_8};
  assign _zz_when_ArraySlice_l173_106_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_107 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_107_1);
  assign _zz_when_ArraySlice_l165_107_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_107_1 = {1'd0, _zz_when_ArraySlice_l165_107_2};
  assign _zz_when_ArraySlice_l166_107 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_107_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_107_2);
  assign _zz_when_ArraySlice_l166_107_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_107_3);
  assign _zz_when_ArraySlice_l166_107_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_107_3 = {1'd0, _zz_when_ArraySlice_l166_107_4};
  assign _zz__zz_when_ArraySlice_l112_107 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_107 = (_zz_when_ArraySlice_l113_107_1 - _zz_when_ArraySlice_l113_107_4);
  assign _zz_when_ArraySlice_l113_107_1 = (_zz_when_ArraySlice_l113_107_2 + _zz_when_ArraySlice_l113_107_3);
  assign _zz_when_ArraySlice_l113_107_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_107_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_107_4 = {1'd0, _zz_when_ArraySlice_l112_107};
  assign _zz__zz_when_ArraySlice_l173_107 = (_zz__zz_when_ArraySlice_l173_107_1 + _zz__zz_when_ArraySlice_l173_107_2);
  assign _zz__zz_when_ArraySlice_l173_107_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_107_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_107_3 = {1'd0, _zz_when_ArraySlice_l112_107};
  assign _zz_when_ArraySlice_l118_107_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_107 = _zz_when_ArraySlice_l118_107_1[5:0];
  assign _zz_when_ArraySlice_l173_107_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_107_1 = {1'd0, _zz_when_ArraySlice_l173_107_2};
  assign _zz_when_ArraySlice_l173_107_3 = (_zz_when_ArraySlice_l173_107_4 + _zz_when_ArraySlice_l173_107_9);
  assign _zz_when_ArraySlice_l173_107_4 = (_zz_when_ArraySlice_l173_107 - _zz_when_ArraySlice_l173_107_5);
  assign _zz_when_ArraySlice_l173_107_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_107_7);
  assign _zz_when_ArraySlice_l173_107_5 = {1'd0, _zz_when_ArraySlice_l173_107_6};
  assign _zz_when_ArraySlice_l173_107_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_107_7 = {1'd0, _zz_when_ArraySlice_l173_107_8};
  assign _zz_when_ArraySlice_l173_107_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_108 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_108_1);
  assign _zz_when_ArraySlice_l165_108_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_108 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_108_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_108_2);
  assign _zz_when_ArraySlice_l166_108_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_108_3);
  assign _zz_when_ArraySlice_l166_108_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_108 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_108 = (_zz_when_ArraySlice_l113_108_1 - _zz_when_ArraySlice_l113_108_4);
  assign _zz_when_ArraySlice_l113_108_1 = (_zz_when_ArraySlice_l113_108_2 + _zz_when_ArraySlice_l113_108_3);
  assign _zz_when_ArraySlice_l113_108_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_108_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_108_4 = {1'd0, _zz_when_ArraySlice_l112_108};
  assign _zz__zz_when_ArraySlice_l173_108 = (_zz__zz_when_ArraySlice_l173_108_1 + _zz__zz_when_ArraySlice_l173_108_2);
  assign _zz__zz_when_ArraySlice_l173_108_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_108_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_108_3 = {1'd0, _zz_when_ArraySlice_l112_108};
  assign _zz_when_ArraySlice_l118_108_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_108 = _zz_when_ArraySlice_l118_108_1[5:0];
  assign _zz_when_ArraySlice_l173_108_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_108_1 = {1'd0, _zz_when_ArraySlice_l173_108_2};
  assign _zz_when_ArraySlice_l173_108_3 = (_zz_when_ArraySlice_l173_108_4 + _zz_when_ArraySlice_l173_108_8);
  assign _zz_when_ArraySlice_l173_108_4 = (_zz_when_ArraySlice_l173_108 - _zz_when_ArraySlice_l173_108_5);
  assign _zz_when_ArraySlice_l173_108_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_108_7);
  assign _zz_when_ArraySlice_l173_108_5 = {1'd0, _zz_when_ArraySlice_l173_108_6};
  assign _zz_when_ArraySlice_l173_108_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_108_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_109 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_109_1);
  assign _zz_when_ArraySlice_l165_109_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_109_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_109 = {1'd0, _zz_when_ArraySlice_l166_109_1};
  assign _zz_when_ArraySlice_l166_109_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_109_3);
  assign _zz_when_ArraySlice_l166_109_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_109_4);
  assign _zz_when_ArraySlice_l166_109_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_109 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_109 = (_zz_when_ArraySlice_l113_109_1 - _zz_when_ArraySlice_l113_109_4);
  assign _zz_when_ArraySlice_l113_109_1 = (_zz_when_ArraySlice_l113_109_2 + _zz_when_ArraySlice_l113_109_3);
  assign _zz_when_ArraySlice_l113_109_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_109_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_109_4 = {1'd0, _zz_when_ArraySlice_l112_109};
  assign _zz__zz_when_ArraySlice_l173_109 = (_zz__zz_when_ArraySlice_l173_109_1 + _zz__zz_when_ArraySlice_l173_109_2);
  assign _zz__zz_when_ArraySlice_l173_109_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_109_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_109_3 = {1'd0, _zz_when_ArraySlice_l112_109};
  assign _zz_when_ArraySlice_l118_109_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_109 = _zz_when_ArraySlice_l118_109_1[5:0];
  assign _zz_when_ArraySlice_l173_109_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_109_1 = {2'd0, _zz_when_ArraySlice_l173_109_2};
  assign _zz_when_ArraySlice_l173_109_3 = (_zz_when_ArraySlice_l173_109_4 + _zz_when_ArraySlice_l173_109_8);
  assign _zz_when_ArraySlice_l173_109_4 = (_zz_when_ArraySlice_l173_109 - _zz_when_ArraySlice_l173_109_5);
  assign _zz_when_ArraySlice_l173_109_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_109_7);
  assign _zz_when_ArraySlice_l173_109_5 = {1'd0, _zz_when_ArraySlice_l173_109_6};
  assign _zz_when_ArraySlice_l173_109_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_109_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_110 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_110_1);
  assign _zz_when_ArraySlice_l165_110_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_110_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_110 = {1'd0, _zz_when_ArraySlice_l166_110_1};
  assign _zz_when_ArraySlice_l166_110_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_110_3);
  assign _zz_when_ArraySlice_l166_110_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_110_4);
  assign _zz_when_ArraySlice_l166_110_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_110 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_110 = (_zz_when_ArraySlice_l113_110_1 - _zz_when_ArraySlice_l113_110_4);
  assign _zz_when_ArraySlice_l113_110_1 = (_zz_when_ArraySlice_l113_110_2 + _zz_when_ArraySlice_l113_110_3);
  assign _zz_when_ArraySlice_l113_110_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_110_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_110_4 = {1'd0, _zz_when_ArraySlice_l112_110};
  assign _zz__zz_when_ArraySlice_l173_110 = (_zz__zz_when_ArraySlice_l173_110_1 + _zz__zz_when_ArraySlice_l173_110_2);
  assign _zz__zz_when_ArraySlice_l173_110_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_110_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_110_3 = {1'd0, _zz_when_ArraySlice_l112_110};
  assign _zz_when_ArraySlice_l118_110_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_110 = _zz_when_ArraySlice_l118_110_1[5:0];
  assign _zz_when_ArraySlice_l173_110_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_110_1 = {2'd0, _zz_when_ArraySlice_l173_110_2};
  assign _zz_when_ArraySlice_l173_110_3 = (_zz_when_ArraySlice_l173_110_4 + _zz_when_ArraySlice_l173_110_8);
  assign _zz_when_ArraySlice_l173_110_4 = (_zz_when_ArraySlice_l173_110 - _zz_when_ArraySlice_l173_110_5);
  assign _zz_when_ArraySlice_l173_110_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_110_7);
  assign _zz_when_ArraySlice_l173_110_5 = {1'd0, _zz_when_ArraySlice_l173_110_6};
  assign _zz_when_ArraySlice_l173_110_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_110_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_111 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_111_1);
  assign _zz_when_ArraySlice_l165_111_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_111_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_111 = {2'd0, _zz_when_ArraySlice_l166_111_1};
  assign _zz_when_ArraySlice_l166_111_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_111_3);
  assign _zz_when_ArraySlice_l166_111_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_111_4);
  assign _zz_when_ArraySlice_l166_111_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_111 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_111 = (_zz_when_ArraySlice_l113_111_1 - _zz_when_ArraySlice_l113_111_4);
  assign _zz_when_ArraySlice_l113_111_1 = (_zz_when_ArraySlice_l113_111_2 + _zz_when_ArraySlice_l113_111_3);
  assign _zz_when_ArraySlice_l113_111_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_111_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_111_4 = {1'd0, _zz_when_ArraySlice_l112_111};
  assign _zz__zz_when_ArraySlice_l173_111 = (_zz__zz_when_ArraySlice_l173_111_1 + _zz__zz_when_ArraySlice_l173_111_2);
  assign _zz__zz_when_ArraySlice_l173_111_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_111_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_111_3 = {1'd0, _zz_when_ArraySlice_l112_111};
  assign _zz_when_ArraySlice_l118_111_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_111 = _zz_when_ArraySlice_l118_111_1[5:0];
  assign _zz_when_ArraySlice_l173_111_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_111_1 = {3'd0, _zz_when_ArraySlice_l173_111_2};
  assign _zz_when_ArraySlice_l173_111_3 = (_zz_when_ArraySlice_l173_111_4 + _zz_when_ArraySlice_l173_111_8);
  assign _zz_when_ArraySlice_l173_111_4 = (_zz_when_ArraySlice_l173_111 - _zz_when_ArraySlice_l173_111_5);
  assign _zz_when_ArraySlice_l173_111_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_111_7);
  assign _zz_when_ArraySlice_l173_111_5 = {1'd0, _zz_when_ArraySlice_l173_111_6};
  assign _zz_when_ArraySlice_l173_111_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_111_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l401_4_1 = (_zz_when_ArraySlice_l401_4_2 + _zz_when_ArraySlice_l401_4_7);
  assign _zz_when_ArraySlice_l401_4_2 = (_zz_when_ArraySlice_l401_4_3 + _zz_when_ArraySlice_l401_4_5);
  assign _zz_when_ArraySlice_l401_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l401_4_4);
  assign _zz_when_ArraySlice_l401_4_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l401_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l401_4_5 = {5'd0, _zz_when_ArraySlice_l401_4_6};
  assign _zz_when_ArraySlice_l401_4_7 = (bReg * 3'b100);
  assign _zz_selectReadFifo_4_15 = 1'b1;
  assign _zz_selectReadFifo_4_14 = {5'd0, _zz_selectReadFifo_4_15};
  assign _zz_when_ArraySlice_l405_4 = (_zz_when_ArraySlice_l405_4_1 % aReg);
  assign _zz_when_ArraySlice_l405_4_1 = (handshakeTimes_4_value + _zz_when_ArraySlice_l405_4_2);
  assign _zz_when_ArraySlice_l405_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l405_4_2 = {12'd0, _zz_when_ArraySlice_l405_4_3};
  assign _zz_when_ArraySlice_l409_4_1 = (selectReadFifo_4 + _zz_when_ArraySlice_l409_4_2);
  assign _zz_when_ArraySlice_l409_4_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l410_4_2 = (_zz_when_ArraySlice_l410_4_3 - _zz_when_ArraySlice_l410_4_4);
  assign _zz_when_ArraySlice_l410_4_1 = {7'd0, _zz_when_ArraySlice_l410_4_2};
  assign _zz_when_ArraySlice_l410_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l410_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l410_4_4 = {5'd0, _zz_when_ArraySlice_l410_4_5};
  assign _zz__zz_when_ArraySlice_l94_13 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_13 = (_zz_when_ArraySlice_l95_13_1 - _zz_when_ArraySlice_l95_13_4);
  assign _zz_when_ArraySlice_l95_13_1 = (_zz_when_ArraySlice_l95_13_2 + _zz_when_ArraySlice_l95_13_3);
  assign _zz_when_ArraySlice_l95_13_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_13_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_13_4 = {1'd0, _zz_when_ArraySlice_l94_13};
  assign _zz__zz_when_ArraySlice_l412_4 = (_zz__zz_when_ArraySlice_l412_4_1 + _zz__zz_when_ArraySlice_l412_4_2);
  assign _zz__zz_when_ArraySlice_l412_4_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l412_4_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l412_4_3 = {1'd0, _zz_when_ArraySlice_l94_13};
  assign _zz_when_ArraySlice_l99_13_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_13 = _zz_when_ArraySlice_l99_13_1[5:0];
  assign _zz_when_ArraySlice_l412_4_1 = (outSliceNumb_4_value + _zz_when_ArraySlice_l412_4_2);
  assign _zz_when_ArraySlice_l412_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l412_4_2 = {6'd0, _zz_when_ArraySlice_l412_4_3};
  assign _zz_when_ArraySlice_l412_4_4 = (_zz_when_ArraySlice_l412_4 / aReg);
  assign _zz_selectReadFifo_4_16 = (selectReadFifo_4 - _zz_selectReadFifo_4_17);
  assign _zz_selectReadFifo_4_17 = {3'd0, bReg};
  assign _zz_selectReadFifo_4_19 = 1'b1;
  assign _zz_selectReadFifo_4_18 = {5'd0, _zz_selectReadFifo_4_19};
  assign _zz_selectReadFifo_4_20 = (selectReadFifo_4 + _zz_selectReadFifo_4_21);
  assign _zz_selectReadFifo_4_21 = (3'b111 * bReg);
  assign _zz_selectReadFifo_4_23 = 1'b1;
  assign _zz_selectReadFifo_4_22 = {5'd0, _zz_selectReadFifo_4_23};
  assign _zz_when_ArraySlice_l165_112 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_112_1);
  assign _zz_when_ArraySlice_l165_112_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_112_1 = {3'd0, _zz_when_ArraySlice_l165_112_2};
  assign _zz_when_ArraySlice_l166_112 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_112_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_112_3);
  assign _zz_when_ArraySlice_l166_112_1 = {1'd0, _zz_when_ArraySlice_l166_112_2};
  assign _zz_when_ArraySlice_l166_112_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_112_4);
  assign _zz_when_ArraySlice_l166_112_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_112_4 = {3'd0, _zz_when_ArraySlice_l166_112_5};
  assign _zz__zz_when_ArraySlice_l112_112 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_112 = (_zz_when_ArraySlice_l113_112_1 - _zz_when_ArraySlice_l113_112_4);
  assign _zz_when_ArraySlice_l113_112_1 = (_zz_when_ArraySlice_l113_112_2 + _zz_when_ArraySlice_l113_112_3);
  assign _zz_when_ArraySlice_l113_112_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_112_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_112_4 = {1'd0, _zz_when_ArraySlice_l112_112};
  assign _zz__zz_when_ArraySlice_l173_112 = (_zz__zz_when_ArraySlice_l173_112_1 + _zz__zz_when_ArraySlice_l173_112_2);
  assign _zz__zz_when_ArraySlice_l173_112_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_112_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_112_3 = {1'd0, _zz_when_ArraySlice_l112_112};
  assign _zz_when_ArraySlice_l118_112_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_112 = _zz_when_ArraySlice_l118_112_1[5:0];
  assign _zz_when_ArraySlice_l173_112_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_112_2 = (_zz_when_ArraySlice_l173_112_3 + _zz_when_ArraySlice_l173_112_8);
  assign _zz_when_ArraySlice_l173_112_3 = (_zz_when_ArraySlice_l173_112 - _zz_when_ArraySlice_l173_112_4);
  assign _zz_when_ArraySlice_l173_112_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_112_6);
  assign _zz_when_ArraySlice_l173_112_4 = {1'd0, _zz_when_ArraySlice_l173_112_5};
  assign _zz_when_ArraySlice_l173_112_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_112_6 = {3'd0, _zz_when_ArraySlice_l173_112_7};
  assign _zz_when_ArraySlice_l173_112_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_113 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_113_1);
  assign _zz_when_ArraySlice_l165_113_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_113_1 = {2'd0, _zz_when_ArraySlice_l165_113_2};
  assign _zz_when_ArraySlice_l166_113 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_113_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_113_2);
  assign _zz_when_ArraySlice_l166_113_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_113_3);
  assign _zz_when_ArraySlice_l166_113_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_113_3 = {2'd0, _zz_when_ArraySlice_l166_113_4};
  assign _zz__zz_when_ArraySlice_l112_113 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_113 = (_zz_when_ArraySlice_l113_113_1 - _zz_when_ArraySlice_l113_113_4);
  assign _zz_when_ArraySlice_l113_113_1 = (_zz_when_ArraySlice_l113_113_2 + _zz_when_ArraySlice_l113_113_3);
  assign _zz_when_ArraySlice_l113_113_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_113_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_113_4 = {1'd0, _zz_when_ArraySlice_l112_113};
  assign _zz__zz_when_ArraySlice_l173_113 = (_zz__zz_when_ArraySlice_l173_113_1 + _zz__zz_when_ArraySlice_l173_113_2);
  assign _zz__zz_when_ArraySlice_l173_113_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_113_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_113_3 = {1'd0, _zz_when_ArraySlice_l112_113};
  assign _zz_when_ArraySlice_l118_113_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_113 = _zz_when_ArraySlice_l118_113_1[5:0];
  assign _zz_when_ArraySlice_l173_113_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_113_1 = {1'd0, _zz_when_ArraySlice_l173_113_2};
  assign _zz_when_ArraySlice_l173_113_3 = (_zz_when_ArraySlice_l173_113_4 + _zz_when_ArraySlice_l173_113_9);
  assign _zz_when_ArraySlice_l173_113_4 = (_zz_when_ArraySlice_l173_113 - _zz_when_ArraySlice_l173_113_5);
  assign _zz_when_ArraySlice_l173_113_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_113_7);
  assign _zz_when_ArraySlice_l173_113_5 = {1'd0, _zz_when_ArraySlice_l173_113_6};
  assign _zz_when_ArraySlice_l173_113_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_113_7 = {2'd0, _zz_when_ArraySlice_l173_113_8};
  assign _zz_when_ArraySlice_l173_113_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_114 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_114_1);
  assign _zz_when_ArraySlice_l165_114_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_114_1 = {1'd0, _zz_when_ArraySlice_l165_114_2};
  assign _zz_when_ArraySlice_l166_114 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_114_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_114_2);
  assign _zz_when_ArraySlice_l166_114_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_114_3);
  assign _zz_when_ArraySlice_l166_114_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_114_3 = {1'd0, _zz_when_ArraySlice_l166_114_4};
  assign _zz__zz_when_ArraySlice_l112_114 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_114 = (_zz_when_ArraySlice_l113_114_1 - _zz_when_ArraySlice_l113_114_4);
  assign _zz_when_ArraySlice_l113_114_1 = (_zz_when_ArraySlice_l113_114_2 + _zz_when_ArraySlice_l113_114_3);
  assign _zz_when_ArraySlice_l113_114_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_114_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_114_4 = {1'd0, _zz_when_ArraySlice_l112_114};
  assign _zz__zz_when_ArraySlice_l173_114 = (_zz__zz_when_ArraySlice_l173_114_1 + _zz__zz_when_ArraySlice_l173_114_2);
  assign _zz__zz_when_ArraySlice_l173_114_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_114_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_114_3 = {1'd0, _zz_when_ArraySlice_l112_114};
  assign _zz_when_ArraySlice_l118_114_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_114 = _zz_when_ArraySlice_l118_114_1[5:0];
  assign _zz_when_ArraySlice_l173_114_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_114_1 = {1'd0, _zz_when_ArraySlice_l173_114_2};
  assign _zz_when_ArraySlice_l173_114_3 = (_zz_when_ArraySlice_l173_114_4 + _zz_when_ArraySlice_l173_114_9);
  assign _zz_when_ArraySlice_l173_114_4 = (_zz_when_ArraySlice_l173_114 - _zz_when_ArraySlice_l173_114_5);
  assign _zz_when_ArraySlice_l173_114_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_114_7);
  assign _zz_when_ArraySlice_l173_114_5 = {1'd0, _zz_when_ArraySlice_l173_114_6};
  assign _zz_when_ArraySlice_l173_114_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_114_7 = {1'd0, _zz_when_ArraySlice_l173_114_8};
  assign _zz_when_ArraySlice_l173_114_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_115 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_115_1);
  assign _zz_when_ArraySlice_l165_115_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_115_1 = {1'd0, _zz_when_ArraySlice_l165_115_2};
  assign _zz_when_ArraySlice_l166_115 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_115_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_115_2);
  assign _zz_when_ArraySlice_l166_115_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_115_3);
  assign _zz_when_ArraySlice_l166_115_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_115_3 = {1'd0, _zz_when_ArraySlice_l166_115_4};
  assign _zz__zz_when_ArraySlice_l112_115 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_115 = (_zz_when_ArraySlice_l113_115_1 - _zz_when_ArraySlice_l113_115_4);
  assign _zz_when_ArraySlice_l113_115_1 = (_zz_when_ArraySlice_l113_115_2 + _zz_when_ArraySlice_l113_115_3);
  assign _zz_when_ArraySlice_l113_115_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_115_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_115_4 = {1'd0, _zz_when_ArraySlice_l112_115};
  assign _zz__zz_when_ArraySlice_l173_115 = (_zz__zz_when_ArraySlice_l173_115_1 + _zz__zz_when_ArraySlice_l173_115_2);
  assign _zz__zz_when_ArraySlice_l173_115_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_115_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_115_3 = {1'd0, _zz_when_ArraySlice_l112_115};
  assign _zz_when_ArraySlice_l118_115_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_115 = _zz_when_ArraySlice_l118_115_1[5:0];
  assign _zz_when_ArraySlice_l173_115_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_115_1 = {1'd0, _zz_when_ArraySlice_l173_115_2};
  assign _zz_when_ArraySlice_l173_115_3 = (_zz_when_ArraySlice_l173_115_4 + _zz_when_ArraySlice_l173_115_9);
  assign _zz_when_ArraySlice_l173_115_4 = (_zz_when_ArraySlice_l173_115 - _zz_when_ArraySlice_l173_115_5);
  assign _zz_when_ArraySlice_l173_115_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_115_7);
  assign _zz_when_ArraySlice_l173_115_5 = {1'd0, _zz_when_ArraySlice_l173_115_6};
  assign _zz_when_ArraySlice_l173_115_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_115_7 = {1'd0, _zz_when_ArraySlice_l173_115_8};
  assign _zz_when_ArraySlice_l173_115_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_116 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_116_1);
  assign _zz_when_ArraySlice_l165_116_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_116 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_116_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_116_2);
  assign _zz_when_ArraySlice_l166_116_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_116_3);
  assign _zz_when_ArraySlice_l166_116_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_116 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_116 = (_zz_when_ArraySlice_l113_116_1 - _zz_when_ArraySlice_l113_116_4);
  assign _zz_when_ArraySlice_l113_116_1 = (_zz_when_ArraySlice_l113_116_2 + _zz_when_ArraySlice_l113_116_3);
  assign _zz_when_ArraySlice_l113_116_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_116_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_116_4 = {1'd0, _zz_when_ArraySlice_l112_116};
  assign _zz__zz_when_ArraySlice_l173_116 = (_zz__zz_when_ArraySlice_l173_116_1 + _zz__zz_when_ArraySlice_l173_116_2);
  assign _zz__zz_when_ArraySlice_l173_116_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_116_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_116_3 = {1'd0, _zz_when_ArraySlice_l112_116};
  assign _zz_when_ArraySlice_l118_116_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_116 = _zz_when_ArraySlice_l118_116_1[5:0];
  assign _zz_when_ArraySlice_l173_116_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_116_1 = {1'd0, _zz_when_ArraySlice_l173_116_2};
  assign _zz_when_ArraySlice_l173_116_3 = (_zz_when_ArraySlice_l173_116_4 + _zz_when_ArraySlice_l173_116_8);
  assign _zz_when_ArraySlice_l173_116_4 = (_zz_when_ArraySlice_l173_116 - _zz_when_ArraySlice_l173_116_5);
  assign _zz_when_ArraySlice_l173_116_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_116_7);
  assign _zz_when_ArraySlice_l173_116_5 = {1'd0, _zz_when_ArraySlice_l173_116_6};
  assign _zz_when_ArraySlice_l173_116_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_116_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_117 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_117_1);
  assign _zz_when_ArraySlice_l165_117_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_117_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_117 = {1'd0, _zz_when_ArraySlice_l166_117_1};
  assign _zz_when_ArraySlice_l166_117_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_117_3);
  assign _zz_when_ArraySlice_l166_117_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_117_4);
  assign _zz_when_ArraySlice_l166_117_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_117 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_117 = (_zz_when_ArraySlice_l113_117_1 - _zz_when_ArraySlice_l113_117_4);
  assign _zz_when_ArraySlice_l113_117_1 = (_zz_when_ArraySlice_l113_117_2 + _zz_when_ArraySlice_l113_117_3);
  assign _zz_when_ArraySlice_l113_117_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_117_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_117_4 = {1'd0, _zz_when_ArraySlice_l112_117};
  assign _zz__zz_when_ArraySlice_l173_117 = (_zz__zz_when_ArraySlice_l173_117_1 + _zz__zz_when_ArraySlice_l173_117_2);
  assign _zz__zz_when_ArraySlice_l173_117_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_117_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_117_3 = {1'd0, _zz_when_ArraySlice_l112_117};
  assign _zz_when_ArraySlice_l118_117_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_117 = _zz_when_ArraySlice_l118_117_1[5:0];
  assign _zz_when_ArraySlice_l173_117_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_117_1 = {2'd0, _zz_when_ArraySlice_l173_117_2};
  assign _zz_when_ArraySlice_l173_117_3 = (_zz_when_ArraySlice_l173_117_4 + _zz_when_ArraySlice_l173_117_8);
  assign _zz_when_ArraySlice_l173_117_4 = (_zz_when_ArraySlice_l173_117 - _zz_when_ArraySlice_l173_117_5);
  assign _zz_when_ArraySlice_l173_117_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_117_7);
  assign _zz_when_ArraySlice_l173_117_5 = {1'd0, _zz_when_ArraySlice_l173_117_6};
  assign _zz_when_ArraySlice_l173_117_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_117_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_118 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_118_1);
  assign _zz_when_ArraySlice_l165_118_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_118_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_118 = {1'd0, _zz_when_ArraySlice_l166_118_1};
  assign _zz_when_ArraySlice_l166_118_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_118_3);
  assign _zz_when_ArraySlice_l166_118_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_118_4);
  assign _zz_when_ArraySlice_l166_118_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_118 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_118 = (_zz_when_ArraySlice_l113_118_1 - _zz_when_ArraySlice_l113_118_4);
  assign _zz_when_ArraySlice_l113_118_1 = (_zz_when_ArraySlice_l113_118_2 + _zz_when_ArraySlice_l113_118_3);
  assign _zz_when_ArraySlice_l113_118_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_118_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_118_4 = {1'd0, _zz_when_ArraySlice_l112_118};
  assign _zz__zz_when_ArraySlice_l173_118 = (_zz__zz_when_ArraySlice_l173_118_1 + _zz__zz_when_ArraySlice_l173_118_2);
  assign _zz__zz_when_ArraySlice_l173_118_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_118_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_118_3 = {1'd0, _zz_when_ArraySlice_l112_118};
  assign _zz_when_ArraySlice_l118_118_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_118 = _zz_when_ArraySlice_l118_118_1[5:0];
  assign _zz_when_ArraySlice_l173_118_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_118_1 = {2'd0, _zz_when_ArraySlice_l173_118_2};
  assign _zz_when_ArraySlice_l173_118_3 = (_zz_when_ArraySlice_l173_118_4 + _zz_when_ArraySlice_l173_118_8);
  assign _zz_when_ArraySlice_l173_118_4 = (_zz_when_ArraySlice_l173_118 - _zz_when_ArraySlice_l173_118_5);
  assign _zz_when_ArraySlice_l173_118_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_118_7);
  assign _zz_when_ArraySlice_l173_118_5 = {1'd0, _zz_when_ArraySlice_l173_118_6};
  assign _zz_when_ArraySlice_l173_118_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_118_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_119 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_119_1);
  assign _zz_when_ArraySlice_l165_119_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_119_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_119 = {2'd0, _zz_when_ArraySlice_l166_119_1};
  assign _zz_when_ArraySlice_l166_119_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_119_3);
  assign _zz_when_ArraySlice_l166_119_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_119_4);
  assign _zz_when_ArraySlice_l166_119_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_119 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_119 = (_zz_when_ArraySlice_l113_119_1 - _zz_when_ArraySlice_l113_119_4);
  assign _zz_when_ArraySlice_l113_119_1 = (_zz_when_ArraySlice_l113_119_2 + _zz_when_ArraySlice_l113_119_3);
  assign _zz_when_ArraySlice_l113_119_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_119_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_119_4 = {1'd0, _zz_when_ArraySlice_l112_119};
  assign _zz__zz_when_ArraySlice_l173_119 = (_zz__zz_when_ArraySlice_l173_119_1 + _zz__zz_when_ArraySlice_l173_119_2);
  assign _zz__zz_when_ArraySlice_l173_119_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_119_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_119_3 = {1'd0, _zz_when_ArraySlice_l112_119};
  assign _zz_when_ArraySlice_l118_119_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_119 = _zz_when_ArraySlice_l118_119_1[5:0];
  assign _zz_when_ArraySlice_l173_119_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_119_1 = {3'd0, _zz_when_ArraySlice_l173_119_2};
  assign _zz_when_ArraySlice_l173_119_3 = (_zz_when_ArraySlice_l173_119_4 + _zz_when_ArraySlice_l173_119_8);
  assign _zz_when_ArraySlice_l173_119_4 = (_zz_when_ArraySlice_l173_119 - _zz_when_ArraySlice_l173_119_5);
  assign _zz_when_ArraySlice_l173_119_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_119_7);
  assign _zz_when_ArraySlice_l173_119_5 = {1'd0, _zz_when_ArraySlice_l173_119_6};
  assign _zz_when_ArraySlice_l173_119_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_119_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l421_4_1 = (_zz_when_ArraySlice_l421_4_2 + _zz_when_ArraySlice_l421_4_7);
  assign _zz_when_ArraySlice_l421_4_2 = (_zz_when_ArraySlice_l421_4_3 + _zz_when_ArraySlice_l421_4_5);
  assign _zz_when_ArraySlice_l421_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l421_4_4);
  assign _zz_when_ArraySlice_l421_4_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l421_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l421_4_5 = {5'd0, _zz_when_ArraySlice_l421_4_6};
  assign _zz_when_ArraySlice_l421_4_7 = (bReg * 3'b100);
  assign _zz_selectReadFifo_4_25 = 1'b1;
  assign _zz_selectReadFifo_4_24 = {5'd0, _zz_selectReadFifo_4_25};
  assign _zz_when_ArraySlice_l425_4 = (_zz_when_ArraySlice_l425_4_1 % aReg);
  assign _zz_when_ArraySlice_l425_4_1 = (handshakeTimes_4_value + _zz_when_ArraySlice_l425_4_2);
  assign _zz_when_ArraySlice_l425_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l425_4_2 = {12'd0, _zz_when_ArraySlice_l425_4_3};
  assign _zz_when_ArraySlice_l436_4_2 = (_zz_when_ArraySlice_l436_4_3 - _zz_when_ArraySlice_l436_4_4);
  assign _zz_when_ArraySlice_l436_4_1 = {7'd0, _zz_when_ArraySlice_l436_4_2};
  assign _zz_when_ArraySlice_l436_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l436_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l436_4_4 = {5'd0, _zz_when_ArraySlice_l436_4_5};
  assign _zz__zz_when_ArraySlice_l94_14 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_14 = (_zz_when_ArraySlice_l95_14_1 - _zz_when_ArraySlice_l95_14_4);
  assign _zz_when_ArraySlice_l95_14_1 = (_zz_when_ArraySlice_l95_14_2 + _zz_when_ArraySlice_l95_14_3);
  assign _zz_when_ArraySlice_l95_14_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_14_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_14_4 = {1'd0, _zz_when_ArraySlice_l94_14};
  assign _zz__zz_when_ArraySlice_l437_4 = (_zz__zz_when_ArraySlice_l437_4_1 + _zz__zz_when_ArraySlice_l437_4_2);
  assign _zz__zz_when_ArraySlice_l437_4_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l437_4_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l437_4_3 = {1'd0, _zz_when_ArraySlice_l94_14};
  assign _zz_when_ArraySlice_l99_14_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_14 = _zz_when_ArraySlice_l99_14_1[5:0];
  assign _zz_when_ArraySlice_l437_4_1 = (outSliceNumb_4_value + _zz_when_ArraySlice_l437_4_2);
  assign _zz_when_ArraySlice_l437_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l437_4_2 = {6'd0, _zz_when_ArraySlice_l437_4_3};
  assign _zz_when_ArraySlice_l437_4_4 = (_zz_when_ArraySlice_l437_4 / aReg);
  assign _zz_selectReadFifo_4_26 = (selectReadFifo_4 - _zz_selectReadFifo_4_27);
  assign _zz_selectReadFifo_4_27 = {3'd0, bReg};
  assign _zz_selectReadFifo_4_29 = 1'b1;
  assign _zz_selectReadFifo_4_28 = {5'd0, _zz_selectReadFifo_4_29};
  assign _zz_when_ArraySlice_l165_120 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_120_1);
  assign _zz_when_ArraySlice_l165_120_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_120_1 = {3'd0, _zz_when_ArraySlice_l165_120_2};
  assign _zz_when_ArraySlice_l166_120 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_120_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_120_3);
  assign _zz_when_ArraySlice_l166_120_1 = {1'd0, _zz_when_ArraySlice_l166_120_2};
  assign _zz_when_ArraySlice_l166_120_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_120_4);
  assign _zz_when_ArraySlice_l166_120_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_120_4 = {3'd0, _zz_when_ArraySlice_l166_120_5};
  assign _zz__zz_when_ArraySlice_l112_120 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_120 = (_zz_when_ArraySlice_l113_120_1 - _zz_when_ArraySlice_l113_120_4);
  assign _zz_when_ArraySlice_l113_120_1 = (_zz_when_ArraySlice_l113_120_2 + _zz_when_ArraySlice_l113_120_3);
  assign _zz_when_ArraySlice_l113_120_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_120_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_120_4 = {1'd0, _zz_when_ArraySlice_l112_120};
  assign _zz__zz_when_ArraySlice_l173_120 = (_zz__zz_when_ArraySlice_l173_120_1 + _zz__zz_when_ArraySlice_l173_120_2);
  assign _zz__zz_when_ArraySlice_l173_120_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_120_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_120_3 = {1'd0, _zz_when_ArraySlice_l112_120};
  assign _zz_when_ArraySlice_l118_120_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_120 = _zz_when_ArraySlice_l118_120_1[5:0];
  assign _zz_when_ArraySlice_l173_120_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_120_2 = (_zz_when_ArraySlice_l173_120_3 + _zz_when_ArraySlice_l173_120_8);
  assign _zz_when_ArraySlice_l173_120_3 = (_zz_when_ArraySlice_l173_120 - _zz_when_ArraySlice_l173_120_4);
  assign _zz_when_ArraySlice_l173_120_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_120_6);
  assign _zz_when_ArraySlice_l173_120_4 = {1'd0, _zz_when_ArraySlice_l173_120_5};
  assign _zz_when_ArraySlice_l173_120_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_120_6 = {3'd0, _zz_when_ArraySlice_l173_120_7};
  assign _zz_when_ArraySlice_l173_120_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_121 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_121_1);
  assign _zz_when_ArraySlice_l165_121_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_121_1 = {2'd0, _zz_when_ArraySlice_l165_121_2};
  assign _zz_when_ArraySlice_l166_121 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_121_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_121_2);
  assign _zz_when_ArraySlice_l166_121_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_121_3);
  assign _zz_when_ArraySlice_l166_121_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_121_3 = {2'd0, _zz_when_ArraySlice_l166_121_4};
  assign _zz__zz_when_ArraySlice_l112_121 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_121 = (_zz_when_ArraySlice_l113_121_1 - _zz_when_ArraySlice_l113_121_4);
  assign _zz_when_ArraySlice_l113_121_1 = (_zz_when_ArraySlice_l113_121_2 + _zz_when_ArraySlice_l113_121_3);
  assign _zz_when_ArraySlice_l113_121_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_121_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_121_4 = {1'd0, _zz_when_ArraySlice_l112_121};
  assign _zz__zz_when_ArraySlice_l173_121 = (_zz__zz_when_ArraySlice_l173_121_1 + _zz__zz_when_ArraySlice_l173_121_2);
  assign _zz__zz_when_ArraySlice_l173_121_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_121_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_121_3 = {1'd0, _zz_when_ArraySlice_l112_121};
  assign _zz_when_ArraySlice_l118_121_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_121 = _zz_when_ArraySlice_l118_121_1[5:0];
  assign _zz_when_ArraySlice_l173_121_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_121_1 = {1'd0, _zz_when_ArraySlice_l173_121_2};
  assign _zz_when_ArraySlice_l173_121_3 = (_zz_when_ArraySlice_l173_121_4 + _zz_when_ArraySlice_l173_121_9);
  assign _zz_when_ArraySlice_l173_121_4 = (_zz_when_ArraySlice_l173_121 - _zz_when_ArraySlice_l173_121_5);
  assign _zz_when_ArraySlice_l173_121_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_121_7);
  assign _zz_when_ArraySlice_l173_121_5 = {1'd0, _zz_when_ArraySlice_l173_121_6};
  assign _zz_when_ArraySlice_l173_121_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_121_7 = {2'd0, _zz_when_ArraySlice_l173_121_8};
  assign _zz_when_ArraySlice_l173_121_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_122 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_122_1);
  assign _zz_when_ArraySlice_l165_122_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_122_1 = {1'd0, _zz_when_ArraySlice_l165_122_2};
  assign _zz_when_ArraySlice_l166_122 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_122_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_122_2);
  assign _zz_when_ArraySlice_l166_122_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_122_3);
  assign _zz_when_ArraySlice_l166_122_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_122_3 = {1'd0, _zz_when_ArraySlice_l166_122_4};
  assign _zz__zz_when_ArraySlice_l112_122 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_122 = (_zz_when_ArraySlice_l113_122_1 - _zz_when_ArraySlice_l113_122_4);
  assign _zz_when_ArraySlice_l113_122_1 = (_zz_when_ArraySlice_l113_122_2 + _zz_when_ArraySlice_l113_122_3);
  assign _zz_when_ArraySlice_l113_122_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_122_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_122_4 = {1'd0, _zz_when_ArraySlice_l112_122};
  assign _zz__zz_when_ArraySlice_l173_122 = (_zz__zz_when_ArraySlice_l173_122_1 + _zz__zz_when_ArraySlice_l173_122_2);
  assign _zz__zz_when_ArraySlice_l173_122_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_122_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_122_3 = {1'd0, _zz_when_ArraySlice_l112_122};
  assign _zz_when_ArraySlice_l118_122_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_122 = _zz_when_ArraySlice_l118_122_1[5:0];
  assign _zz_when_ArraySlice_l173_122_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_122_1 = {1'd0, _zz_when_ArraySlice_l173_122_2};
  assign _zz_when_ArraySlice_l173_122_3 = (_zz_when_ArraySlice_l173_122_4 + _zz_when_ArraySlice_l173_122_9);
  assign _zz_when_ArraySlice_l173_122_4 = (_zz_when_ArraySlice_l173_122 - _zz_when_ArraySlice_l173_122_5);
  assign _zz_when_ArraySlice_l173_122_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_122_7);
  assign _zz_when_ArraySlice_l173_122_5 = {1'd0, _zz_when_ArraySlice_l173_122_6};
  assign _zz_when_ArraySlice_l173_122_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_122_7 = {1'd0, _zz_when_ArraySlice_l173_122_8};
  assign _zz_when_ArraySlice_l173_122_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_123 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_123_1);
  assign _zz_when_ArraySlice_l165_123_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_123_1 = {1'd0, _zz_when_ArraySlice_l165_123_2};
  assign _zz_when_ArraySlice_l166_123 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_123_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_123_2);
  assign _zz_when_ArraySlice_l166_123_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_123_3);
  assign _zz_when_ArraySlice_l166_123_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_123_3 = {1'd0, _zz_when_ArraySlice_l166_123_4};
  assign _zz__zz_when_ArraySlice_l112_123 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_123 = (_zz_when_ArraySlice_l113_123_1 - _zz_when_ArraySlice_l113_123_4);
  assign _zz_when_ArraySlice_l113_123_1 = (_zz_when_ArraySlice_l113_123_2 + _zz_when_ArraySlice_l113_123_3);
  assign _zz_when_ArraySlice_l113_123_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_123_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_123_4 = {1'd0, _zz_when_ArraySlice_l112_123};
  assign _zz__zz_when_ArraySlice_l173_123 = (_zz__zz_when_ArraySlice_l173_123_1 + _zz__zz_when_ArraySlice_l173_123_2);
  assign _zz__zz_when_ArraySlice_l173_123_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_123_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_123_3 = {1'd0, _zz_when_ArraySlice_l112_123};
  assign _zz_when_ArraySlice_l118_123_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_123 = _zz_when_ArraySlice_l118_123_1[5:0];
  assign _zz_when_ArraySlice_l173_123_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_123_1 = {1'd0, _zz_when_ArraySlice_l173_123_2};
  assign _zz_when_ArraySlice_l173_123_3 = (_zz_when_ArraySlice_l173_123_4 + _zz_when_ArraySlice_l173_123_9);
  assign _zz_when_ArraySlice_l173_123_4 = (_zz_when_ArraySlice_l173_123 - _zz_when_ArraySlice_l173_123_5);
  assign _zz_when_ArraySlice_l173_123_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_123_7);
  assign _zz_when_ArraySlice_l173_123_5 = {1'd0, _zz_when_ArraySlice_l173_123_6};
  assign _zz_when_ArraySlice_l173_123_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_123_7 = {1'd0, _zz_when_ArraySlice_l173_123_8};
  assign _zz_when_ArraySlice_l173_123_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_124 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_124_1);
  assign _zz_when_ArraySlice_l165_124_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_124 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_124_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_124_2);
  assign _zz_when_ArraySlice_l166_124_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_124_3);
  assign _zz_when_ArraySlice_l166_124_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_124 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_124 = (_zz_when_ArraySlice_l113_124_1 - _zz_when_ArraySlice_l113_124_4);
  assign _zz_when_ArraySlice_l113_124_1 = (_zz_when_ArraySlice_l113_124_2 + _zz_when_ArraySlice_l113_124_3);
  assign _zz_when_ArraySlice_l113_124_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_124_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_124_4 = {1'd0, _zz_when_ArraySlice_l112_124};
  assign _zz__zz_when_ArraySlice_l173_124 = (_zz__zz_when_ArraySlice_l173_124_1 + _zz__zz_when_ArraySlice_l173_124_2);
  assign _zz__zz_when_ArraySlice_l173_124_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_124_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_124_3 = {1'd0, _zz_when_ArraySlice_l112_124};
  assign _zz_when_ArraySlice_l118_124_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_124 = _zz_when_ArraySlice_l118_124_1[5:0];
  assign _zz_when_ArraySlice_l173_124_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_124_1 = {1'd0, _zz_when_ArraySlice_l173_124_2};
  assign _zz_when_ArraySlice_l173_124_3 = (_zz_when_ArraySlice_l173_124_4 + _zz_when_ArraySlice_l173_124_8);
  assign _zz_when_ArraySlice_l173_124_4 = (_zz_when_ArraySlice_l173_124 - _zz_when_ArraySlice_l173_124_5);
  assign _zz_when_ArraySlice_l173_124_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_124_7);
  assign _zz_when_ArraySlice_l173_124_5 = {1'd0, _zz_when_ArraySlice_l173_124_6};
  assign _zz_when_ArraySlice_l173_124_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_124_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_125 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_125_1);
  assign _zz_when_ArraySlice_l165_125_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_125_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_125 = {1'd0, _zz_when_ArraySlice_l166_125_1};
  assign _zz_when_ArraySlice_l166_125_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_125_3);
  assign _zz_when_ArraySlice_l166_125_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_125_4);
  assign _zz_when_ArraySlice_l166_125_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_125 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_125 = (_zz_when_ArraySlice_l113_125_1 - _zz_when_ArraySlice_l113_125_4);
  assign _zz_when_ArraySlice_l113_125_1 = (_zz_when_ArraySlice_l113_125_2 + _zz_when_ArraySlice_l113_125_3);
  assign _zz_when_ArraySlice_l113_125_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_125_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_125_4 = {1'd0, _zz_when_ArraySlice_l112_125};
  assign _zz__zz_when_ArraySlice_l173_125 = (_zz__zz_when_ArraySlice_l173_125_1 + _zz__zz_when_ArraySlice_l173_125_2);
  assign _zz__zz_when_ArraySlice_l173_125_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_125_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_125_3 = {1'd0, _zz_when_ArraySlice_l112_125};
  assign _zz_when_ArraySlice_l118_125_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_125 = _zz_when_ArraySlice_l118_125_1[5:0];
  assign _zz_when_ArraySlice_l173_125_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_125_1 = {2'd0, _zz_when_ArraySlice_l173_125_2};
  assign _zz_when_ArraySlice_l173_125_3 = (_zz_when_ArraySlice_l173_125_4 + _zz_when_ArraySlice_l173_125_8);
  assign _zz_when_ArraySlice_l173_125_4 = (_zz_when_ArraySlice_l173_125 - _zz_when_ArraySlice_l173_125_5);
  assign _zz_when_ArraySlice_l173_125_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_125_7);
  assign _zz_when_ArraySlice_l173_125_5 = {1'd0, _zz_when_ArraySlice_l173_125_6};
  assign _zz_when_ArraySlice_l173_125_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_125_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_126 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_126_1);
  assign _zz_when_ArraySlice_l165_126_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_126_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_126 = {1'd0, _zz_when_ArraySlice_l166_126_1};
  assign _zz_when_ArraySlice_l166_126_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_126_3);
  assign _zz_when_ArraySlice_l166_126_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_126_4);
  assign _zz_when_ArraySlice_l166_126_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_126 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_126 = (_zz_when_ArraySlice_l113_126_1 - _zz_when_ArraySlice_l113_126_4);
  assign _zz_when_ArraySlice_l113_126_1 = (_zz_when_ArraySlice_l113_126_2 + _zz_when_ArraySlice_l113_126_3);
  assign _zz_when_ArraySlice_l113_126_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_126_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_126_4 = {1'd0, _zz_when_ArraySlice_l112_126};
  assign _zz__zz_when_ArraySlice_l173_126 = (_zz__zz_when_ArraySlice_l173_126_1 + _zz__zz_when_ArraySlice_l173_126_2);
  assign _zz__zz_when_ArraySlice_l173_126_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_126_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_126_3 = {1'd0, _zz_when_ArraySlice_l112_126};
  assign _zz_when_ArraySlice_l118_126_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_126 = _zz_when_ArraySlice_l118_126_1[5:0];
  assign _zz_when_ArraySlice_l173_126_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_126_1 = {2'd0, _zz_when_ArraySlice_l173_126_2};
  assign _zz_when_ArraySlice_l173_126_3 = (_zz_when_ArraySlice_l173_126_4 + _zz_when_ArraySlice_l173_126_8);
  assign _zz_when_ArraySlice_l173_126_4 = (_zz_when_ArraySlice_l173_126 - _zz_when_ArraySlice_l173_126_5);
  assign _zz_when_ArraySlice_l173_126_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_126_7);
  assign _zz_when_ArraySlice_l173_126_5 = {1'd0, _zz_when_ArraySlice_l173_126_6};
  assign _zz_when_ArraySlice_l173_126_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_126_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_127 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_127_1);
  assign _zz_when_ArraySlice_l165_127_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_127_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_127 = {2'd0, _zz_when_ArraySlice_l166_127_1};
  assign _zz_when_ArraySlice_l166_127_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_127_3);
  assign _zz_when_ArraySlice_l166_127_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_127_4);
  assign _zz_when_ArraySlice_l166_127_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_127 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_127 = (_zz_when_ArraySlice_l113_127_1 - _zz_when_ArraySlice_l113_127_4);
  assign _zz_when_ArraySlice_l113_127_1 = (_zz_when_ArraySlice_l113_127_2 + _zz_when_ArraySlice_l113_127_3);
  assign _zz_when_ArraySlice_l113_127_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_127_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_127_4 = {1'd0, _zz_when_ArraySlice_l112_127};
  assign _zz__zz_when_ArraySlice_l173_127 = (_zz__zz_when_ArraySlice_l173_127_1 + _zz__zz_when_ArraySlice_l173_127_2);
  assign _zz__zz_when_ArraySlice_l173_127_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_127_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_127_3 = {1'd0, _zz_when_ArraySlice_l112_127};
  assign _zz_when_ArraySlice_l118_127_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_127 = _zz_when_ArraySlice_l118_127_1[5:0];
  assign _zz_when_ArraySlice_l173_127_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_127_1 = {3'd0, _zz_when_ArraySlice_l173_127_2};
  assign _zz_when_ArraySlice_l173_127_3 = (_zz_when_ArraySlice_l173_127_4 + _zz_when_ArraySlice_l173_127_8);
  assign _zz_when_ArraySlice_l173_127_4 = (_zz_when_ArraySlice_l173_127 - _zz_when_ArraySlice_l173_127_5);
  assign _zz_when_ArraySlice_l173_127_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_127_7);
  assign _zz_when_ArraySlice_l173_127_5 = {1'd0, _zz_when_ArraySlice_l173_127_6};
  assign _zz_when_ArraySlice_l173_127_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_127_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_4_31 = 1'b1;
  assign _zz_selectReadFifo_4_30 = {5'd0, _zz_selectReadFifo_4_31};
  assign _zz_when_ArraySlice_l448_4 = (_zz_when_ArraySlice_l448_4_1 % aReg);
  assign _zz_when_ArraySlice_l448_4_1 = (handshakeTimes_4_value + _zz_when_ArraySlice_l448_4_2);
  assign _zz_when_ArraySlice_l448_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l448_4_2 = {12'd0, _zz_when_ArraySlice_l448_4_3};
  assign _zz_when_ArraySlice_l434_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l434_4_1);
  assign _zz_when_ArraySlice_l434_4_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l455_4_2 = (_zz_when_ArraySlice_l455_4_3 - _zz_when_ArraySlice_l455_4_4);
  assign _zz_when_ArraySlice_l455_4_1 = {7'd0, _zz_when_ArraySlice_l455_4_2};
  assign _zz_when_ArraySlice_l455_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l455_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l455_4_4 = {5'd0, _zz_when_ArraySlice_l455_4_5};
  assign _zz_when_ArraySlice_l373_5 = (selectReadFifo_5 + _zz_when_ArraySlice_l373_5_1);
  assign _zz_when_ArraySlice_l373_5_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l374_5_1 = (selectReadFifo_5 + _zz_when_ArraySlice_l374_5_2);
  assign _zz_when_ArraySlice_l374_5_2 = (bReg * 3'b101);
  assign _zz__zz_outputStreamArrayData_5_valid = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l380_5_2 = 1'b1;
  assign _zz_when_ArraySlice_l380_5_1 = {6'd0, _zz_when_ArraySlice_l380_5_2};
  assign _zz_when_ArraySlice_l380_5_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l380_5_5);
  assign _zz_when_ArraySlice_l380_5_5 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l381_5_1 = (_zz_when_ArraySlice_l381_5_2 - _zz_when_ArraySlice_l381_5_3);
  assign _zz_when_ArraySlice_l381_5 = {7'd0, _zz_when_ArraySlice_l381_5_1};
  assign _zz_when_ArraySlice_l381_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l381_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l381_5_3 = {5'd0, _zz_when_ArraySlice_l381_5_4};
  assign _zz_selectReadFifo_5 = (selectReadFifo_5 - _zz_selectReadFifo_5_1);
  assign _zz_selectReadFifo_5_1 = {3'd0, bReg};
  assign _zz_selectReadFifo_5_3 = 1'b1;
  assign _zz_selectReadFifo_5_2 = {5'd0, _zz_selectReadFifo_5_3};
  assign _zz_selectReadFifo_5_5 = 1'b1;
  assign _zz_selectReadFifo_5_4 = {5'd0, _zz_selectReadFifo_5_5};
  assign _zz_when_ArraySlice_l384_5 = (_zz_when_ArraySlice_l384_5_1 % aReg);
  assign _zz_when_ArraySlice_l384_5_1 = (handshakeTimes_5_value + _zz_when_ArraySlice_l384_5_2);
  assign _zz_when_ArraySlice_l384_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l384_5_2 = {12'd0, _zz_when_ArraySlice_l384_5_3};
  assign _zz_when_ArraySlice_l389_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l389_5_3);
  assign _zz_when_ArraySlice_l389_5_3 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l389_5_5 = 1'b1;
  assign _zz_when_ArraySlice_l389_5_4 = {6'd0, _zz_when_ArraySlice_l389_5_5};
  assign _zz_when_ArraySlice_l390_5_1 = (_zz_when_ArraySlice_l390_5_2 - _zz_when_ArraySlice_l390_5_3);
  assign _zz_when_ArraySlice_l390_5 = {7'd0, _zz_when_ArraySlice_l390_5_1};
  assign _zz_when_ArraySlice_l390_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l390_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l390_5_3 = {5'd0, _zz_when_ArraySlice_l390_5_4};
  assign _zz__zz_when_ArraySlice_l94_15 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_15 = (_zz_when_ArraySlice_l95_15_1 - _zz_when_ArraySlice_l95_15_4);
  assign _zz_when_ArraySlice_l95_15_1 = (_zz_when_ArraySlice_l95_15_2 + _zz_when_ArraySlice_l95_15_3);
  assign _zz_when_ArraySlice_l95_15_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_15_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_15_4 = {1'd0, _zz_when_ArraySlice_l94_15};
  assign _zz__zz_when_ArraySlice_l392_5 = (_zz__zz_when_ArraySlice_l392_5_1 + _zz__zz_when_ArraySlice_l392_5_2);
  assign _zz__zz_when_ArraySlice_l392_5_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l392_5_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l392_5_3 = {1'd0, _zz_when_ArraySlice_l94_15};
  assign _zz_when_ArraySlice_l99_15_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_15 = _zz_when_ArraySlice_l99_15_1[5:0];
  assign _zz_when_ArraySlice_l392_5_1 = (outSliceNumb_5_value + _zz_when_ArraySlice_l392_5_2);
  assign _zz_when_ArraySlice_l392_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l392_5_2 = {6'd0, _zz_when_ArraySlice_l392_5_3};
  assign _zz_when_ArraySlice_l392_5_4 = (_zz_when_ArraySlice_l392_5 / aReg);
  assign _zz_selectReadFifo_5_6 = (selectReadFifo_5 - _zz_selectReadFifo_5_7);
  assign _zz_selectReadFifo_5_7 = {3'd0, bReg};
  assign _zz_selectReadFifo_5_9 = 1'b1;
  assign _zz_selectReadFifo_5_8 = {5'd0, _zz_selectReadFifo_5_9};
  assign _zz_selectReadFifo_5_10 = (selectReadFifo_5 + _zz_selectReadFifo_5_11);
  assign _zz_selectReadFifo_5_11 = (3'b111 * bReg);
  assign _zz_selectReadFifo_5_13 = 1'b1;
  assign _zz_selectReadFifo_5_12 = {5'd0, _zz_selectReadFifo_5_13};
  assign _zz_when_ArraySlice_l165_128 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_128_1);
  assign _zz_when_ArraySlice_l165_128_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_128_1 = {3'd0, _zz_when_ArraySlice_l165_128_2};
  assign _zz_when_ArraySlice_l166_128 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_128_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_128_3);
  assign _zz_when_ArraySlice_l166_128_1 = {1'd0, _zz_when_ArraySlice_l166_128_2};
  assign _zz_when_ArraySlice_l166_128_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_128_4);
  assign _zz_when_ArraySlice_l166_128_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_128_4 = {3'd0, _zz_when_ArraySlice_l166_128_5};
  assign _zz__zz_when_ArraySlice_l112_128 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_128 = (_zz_when_ArraySlice_l113_128_1 - _zz_when_ArraySlice_l113_128_4);
  assign _zz_when_ArraySlice_l113_128_1 = (_zz_when_ArraySlice_l113_128_2 + _zz_when_ArraySlice_l113_128_3);
  assign _zz_when_ArraySlice_l113_128_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_128_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_128_4 = {1'd0, _zz_when_ArraySlice_l112_128};
  assign _zz__zz_when_ArraySlice_l173_128 = (_zz__zz_when_ArraySlice_l173_128_1 + _zz__zz_when_ArraySlice_l173_128_2);
  assign _zz__zz_when_ArraySlice_l173_128_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_128_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_128_3 = {1'd0, _zz_when_ArraySlice_l112_128};
  assign _zz_when_ArraySlice_l118_128_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_128 = _zz_when_ArraySlice_l118_128_1[5:0];
  assign _zz_when_ArraySlice_l173_128_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_128_2 = (_zz_when_ArraySlice_l173_128_3 + _zz_when_ArraySlice_l173_128_8);
  assign _zz_when_ArraySlice_l173_128_3 = (_zz_when_ArraySlice_l173_128 - _zz_when_ArraySlice_l173_128_4);
  assign _zz_when_ArraySlice_l173_128_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_128_6);
  assign _zz_when_ArraySlice_l173_128_4 = {1'd0, _zz_when_ArraySlice_l173_128_5};
  assign _zz_when_ArraySlice_l173_128_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_128_6 = {3'd0, _zz_when_ArraySlice_l173_128_7};
  assign _zz_when_ArraySlice_l173_128_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_129 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_129_1);
  assign _zz_when_ArraySlice_l165_129_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_129_1 = {2'd0, _zz_when_ArraySlice_l165_129_2};
  assign _zz_when_ArraySlice_l166_129 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_129_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_129_2);
  assign _zz_when_ArraySlice_l166_129_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_129_3);
  assign _zz_when_ArraySlice_l166_129_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_129_3 = {2'd0, _zz_when_ArraySlice_l166_129_4};
  assign _zz__zz_when_ArraySlice_l112_129 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_129 = (_zz_when_ArraySlice_l113_129_1 - _zz_when_ArraySlice_l113_129_4);
  assign _zz_when_ArraySlice_l113_129_1 = (_zz_when_ArraySlice_l113_129_2 + _zz_when_ArraySlice_l113_129_3);
  assign _zz_when_ArraySlice_l113_129_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_129_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_129_4 = {1'd0, _zz_when_ArraySlice_l112_129};
  assign _zz__zz_when_ArraySlice_l173_129 = (_zz__zz_when_ArraySlice_l173_129_1 + _zz__zz_when_ArraySlice_l173_129_2);
  assign _zz__zz_when_ArraySlice_l173_129_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_129_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_129_3 = {1'd0, _zz_when_ArraySlice_l112_129};
  assign _zz_when_ArraySlice_l118_129_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_129 = _zz_when_ArraySlice_l118_129_1[5:0];
  assign _zz_when_ArraySlice_l173_129_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_129_1 = {1'd0, _zz_when_ArraySlice_l173_129_2};
  assign _zz_when_ArraySlice_l173_129_3 = (_zz_when_ArraySlice_l173_129_4 + _zz_when_ArraySlice_l173_129_9);
  assign _zz_when_ArraySlice_l173_129_4 = (_zz_when_ArraySlice_l173_129 - _zz_when_ArraySlice_l173_129_5);
  assign _zz_when_ArraySlice_l173_129_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_129_7);
  assign _zz_when_ArraySlice_l173_129_5 = {1'd0, _zz_when_ArraySlice_l173_129_6};
  assign _zz_when_ArraySlice_l173_129_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_129_7 = {2'd0, _zz_when_ArraySlice_l173_129_8};
  assign _zz_when_ArraySlice_l173_129_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_130 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_130_1);
  assign _zz_when_ArraySlice_l165_130_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_130_1 = {1'd0, _zz_when_ArraySlice_l165_130_2};
  assign _zz_when_ArraySlice_l166_130 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_130_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_130_2);
  assign _zz_when_ArraySlice_l166_130_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_130_3);
  assign _zz_when_ArraySlice_l166_130_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_130_3 = {1'd0, _zz_when_ArraySlice_l166_130_4};
  assign _zz__zz_when_ArraySlice_l112_130 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_130 = (_zz_when_ArraySlice_l113_130_1 - _zz_when_ArraySlice_l113_130_4);
  assign _zz_when_ArraySlice_l113_130_1 = (_zz_when_ArraySlice_l113_130_2 + _zz_when_ArraySlice_l113_130_3);
  assign _zz_when_ArraySlice_l113_130_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_130_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_130_4 = {1'd0, _zz_when_ArraySlice_l112_130};
  assign _zz__zz_when_ArraySlice_l173_130 = (_zz__zz_when_ArraySlice_l173_130_1 + _zz__zz_when_ArraySlice_l173_130_2);
  assign _zz__zz_when_ArraySlice_l173_130_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_130_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_130_3 = {1'd0, _zz_when_ArraySlice_l112_130};
  assign _zz_when_ArraySlice_l118_130_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_130 = _zz_when_ArraySlice_l118_130_1[5:0];
  assign _zz_when_ArraySlice_l173_130_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_130_1 = {1'd0, _zz_when_ArraySlice_l173_130_2};
  assign _zz_when_ArraySlice_l173_130_3 = (_zz_when_ArraySlice_l173_130_4 + _zz_when_ArraySlice_l173_130_9);
  assign _zz_when_ArraySlice_l173_130_4 = (_zz_when_ArraySlice_l173_130 - _zz_when_ArraySlice_l173_130_5);
  assign _zz_when_ArraySlice_l173_130_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_130_7);
  assign _zz_when_ArraySlice_l173_130_5 = {1'd0, _zz_when_ArraySlice_l173_130_6};
  assign _zz_when_ArraySlice_l173_130_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_130_7 = {1'd0, _zz_when_ArraySlice_l173_130_8};
  assign _zz_when_ArraySlice_l173_130_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_131 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_131_1);
  assign _zz_when_ArraySlice_l165_131_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_131_1 = {1'd0, _zz_when_ArraySlice_l165_131_2};
  assign _zz_when_ArraySlice_l166_131 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_131_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_131_2);
  assign _zz_when_ArraySlice_l166_131_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_131_3);
  assign _zz_when_ArraySlice_l166_131_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_131_3 = {1'd0, _zz_when_ArraySlice_l166_131_4};
  assign _zz__zz_when_ArraySlice_l112_131 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_131 = (_zz_when_ArraySlice_l113_131_1 - _zz_when_ArraySlice_l113_131_4);
  assign _zz_when_ArraySlice_l113_131_1 = (_zz_when_ArraySlice_l113_131_2 + _zz_when_ArraySlice_l113_131_3);
  assign _zz_when_ArraySlice_l113_131_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_131_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_131_4 = {1'd0, _zz_when_ArraySlice_l112_131};
  assign _zz__zz_when_ArraySlice_l173_131 = (_zz__zz_when_ArraySlice_l173_131_1 + _zz__zz_when_ArraySlice_l173_131_2);
  assign _zz__zz_when_ArraySlice_l173_131_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_131_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_131_3 = {1'd0, _zz_when_ArraySlice_l112_131};
  assign _zz_when_ArraySlice_l118_131_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_131 = _zz_when_ArraySlice_l118_131_1[5:0];
  assign _zz_when_ArraySlice_l173_131_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_131_1 = {1'd0, _zz_when_ArraySlice_l173_131_2};
  assign _zz_when_ArraySlice_l173_131_3 = (_zz_when_ArraySlice_l173_131_4 + _zz_when_ArraySlice_l173_131_9);
  assign _zz_when_ArraySlice_l173_131_4 = (_zz_when_ArraySlice_l173_131 - _zz_when_ArraySlice_l173_131_5);
  assign _zz_when_ArraySlice_l173_131_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_131_7);
  assign _zz_when_ArraySlice_l173_131_5 = {1'd0, _zz_when_ArraySlice_l173_131_6};
  assign _zz_when_ArraySlice_l173_131_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_131_7 = {1'd0, _zz_when_ArraySlice_l173_131_8};
  assign _zz_when_ArraySlice_l173_131_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_132 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_132_1);
  assign _zz_when_ArraySlice_l165_132_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_132 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_132_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_132_2);
  assign _zz_when_ArraySlice_l166_132_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_132_3);
  assign _zz_when_ArraySlice_l166_132_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_132 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_132 = (_zz_when_ArraySlice_l113_132_1 - _zz_when_ArraySlice_l113_132_4);
  assign _zz_when_ArraySlice_l113_132_1 = (_zz_when_ArraySlice_l113_132_2 + _zz_when_ArraySlice_l113_132_3);
  assign _zz_when_ArraySlice_l113_132_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_132_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_132_4 = {1'd0, _zz_when_ArraySlice_l112_132};
  assign _zz__zz_when_ArraySlice_l173_132 = (_zz__zz_when_ArraySlice_l173_132_1 + _zz__zz_when_ArraySlice_l173_132_2);
  assign _zz__zz_when_ArraySlice_l173_132_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_132_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_132_3 = {1'd0, _zz_when_ArraySlice_l112_132};
  assign _zz_when_ArraySlice_l118_132_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_132 = _zz_when_ArraySlice_l118_132_1[5:0];
  assign _zz_when_ArraySlice_l173_132_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_132_1 = {1'd0, _zz_when_ArraySlice_l173_132_2};
  assign _zz_when_ArraySlice_l173_132_3 = (_zz_when_ArraySlice_l173_132_4 + _zz_when_ArraySlice_l173_132_8);
  assign _zz_when_ArraySlice_l173_132_4 = (_zz_when_ArraySlice_l173_132 - _zz_when_ArraySlice_l173_132_5);
  assign _zz_when_ArraySlice_l173_132_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_132_7);
  assign _zz_when_ArraySlice_l173_132_5 = {1'd0, _zz_when_ArraySlice_l173_132_6};
  assign _zz_when_ArraySlice_l173_132_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_132_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_133 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_133_1);
  assign _zz_when_ArraySlice_l165_133_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_133_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_133 = {1'd0, _zz_when_ArraySlice_l166_133_1};
  assign _zz_when_ArraySlice_l166_133_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_133_3);
  assign _zz_when_ArraySlice_l166_133_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_133_4);
  assign _zz_when_ArraySlice_l166_133_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_133 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_133 = (_zz_when_ArraySlice_l113_133_1 - _zz_when_ArraySlice_l113_133_4);
  assign _zz_when_ArraySlice_l113_133_1 = (_zz_when_ArraySlice_l113_133_2 + _zz_when_ArraySlice_l113_133_3);
  assign _zz_when_ArraySlice_l113_133_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_133_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_133_4 = {1'd0, _zz_when_ArraySlice_l112_133};
  assign _zz__zz_when_ArraySlice_l173_133 = (_zz__zz_when_ArraySlice_l173_133_1 + _zz__zz_when_ArraySlice_l173_133_2);
  assign _zz__zz_when_ArraySlice_l173_133_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_133_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_133_3 = {1'd0, _zz_when_ArraySlice_l112_133};
  assign _zz_when_ArraySlice_l118_133_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_133 = _zz_when_ArraySlice_l118_133_1[5:0];
  assign _zz_when_ArraySlice_l173_133_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_133_1 = {2'd0, _zz_when_ArraySlice_l173_133_2};
  assign _zz_when_ArraySlice_l173_133_3 = (_zz_when_ArraySlice_l173_133_4 + _zz_when_ArraySlice_l173_133_8);
  assign _zz_when_ArraySlice_l173_133_4 = (_zz_when_ArraySlice_l173_133 - _zz_when_ArraySlice_l173_133_5);
  assign _zz_when_ArraySlice_l173_133_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_133_7);
  assign _zz_when_ArraySlice_l173_133_5 = {1'd0, _zz_when_ArraySlice_l173_133_6};
  assign _zz_when_ArraySlice_l173_133_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_133_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_134 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_134_1);
  assign _zz_when_ArraySlice_l165_134_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_134_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_134 = {1'd0, _zz_when_ArraySlice_l166_134_1};
  assign _zz_when_ArraySlice_l166_134_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_134_3);
  assign _zz_when_ArraySlice_l166_134_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_134_4);
  assign _zz_when_ArraySlice_l166_134_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_134 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_134 = (_zz_when_ArraySlice_l113_134_1 - _zz_when_ArraySlice_l113_134_4);
  assign _zz_when_ArraySlice_l113_134_1 = (_zz_when_ArraySlice_l113_134_2 + _zz_when_ArraySlice_l113_134_3);
  assign _zz_when_ArraySlice_l113_134_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_134_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_134_4 = {1'd0, _zz_when_ArraySlice_l112_134};
  assign _zz__zz_when_ArraySlice_l173_134 = (_zz__zz_when_ArraySlice_l173_134_1 + _zz__zz_when_ArraySlice_l173_134_2);
  assign _zz__zz_when_ArraySlice_l173_134_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_134_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_134_3 = {1'd0, _zz_when_ArraySlice_l112_134};
  assign _zz_when_ArraySlice_l118_134_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_134 = _zz_when_ArraySlice_l118_134_1[5:0];
  assign _zz_when_ArraySlice_l173_134_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_134_1 = {2'd0, _zz_when_ArraySlice_l173_134_2};
  assign _zz_when_ArraySlice_l173_134_3 = (_zz_when_ArraySlice_l173_134_4 + _zz_when_ArraySlice_l173_134_8);
  assign _zz_when_ArraySlice_l173_134_4 = (_zz_when_ArraySlice_l173_134 - _zz_when_ArraySlice_l173_134_5);
  assign _zz_when_ArraySlice_l173_134_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_134_7);
  assign _zz_when_ArraySlice_l173_134_5 = {1'd0, _zz_when_ArraySlice_l173_134_6};
  assign _zz_when_ArraySlice_l173_134_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_134_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_135 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_135_1);
  assign _zz_when_ArraySlice_l165_135_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_135_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_135 = {2'd0, _zz_when_ArraySlice_l166_135_1};
  assign _zz_when_ArraySlice_l166_135_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_135_3);
  assign _zz_when_ArraySlice_l166_135_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_135_4);
  assign _zz_when_ArraySlice_l166_135_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_135 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_135 = (_zz_when_ArraySlice_l113_135_1 - _zz_when_ArraySlice_l113_135_4);
  assign _zz_when_ArraySlice_l113_135_1 = (_zz_when_ArraySlice_l113_135_2 + _zz_when_ArraySlice_l113_135_3);
  assign _zz_when_ArraySlice_l113_135_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_135_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_135_4 = {1'd0, _zz_when_ArraySlice_l112_135};
  assign _zz__zz_when_ArraySlice_l173_135 = (_zz__zz_when_ArraySlice_l173_135_1 + _zz__zz_when_ArraySlice_l173_135_2);
  assign _zz__zz_when_ArraySlice_l173_135_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_135_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_135_3 = {1'd0, _zz_when_ArraySlice_l112_135};
  assign _zz_when_ArraySlice_l118_135_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_135 = _zz_when_ArraySlice_l118_135_1[5:0];
  assign _zz_when_ArraySlice_l173_135_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_135_1 = {3'd0, _zz_when_ArraySlice_l173_135_2};
  assign _zz_when_ArraySlice_l173_135_3 = (_zz_when_ArraySlice_l173_135_4 + _zz_when_ArraySlice_l173_135_8);
  assign _zz_when_ArraySlice_l173_135_4 = (_zz_when_ArraySlice_l173_135 - _zz_when_ArraySlice_l173_135_5);
  assign _zz_when_ArraySlice_l173_135_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_135_7);
  assign _zz_when_ArraySlice_l173_135_5 = {1'd0, _zz_when_ArraySlice_l173_135_6};
  assign _zz_when_ArraySlice_l173_135_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_135_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l401_5_1 = (_zz_when_ArraySlice_l401_5_2 + _zz_when_ArraySlice_l401_5_7);
  assign _zz_when_ArraySlice_l401_5_2 = (_zz_when_ArraySlice_l401_5_3 + _zz_when_ArraySlice_l401_5_5);
  assign _zz_when_ArraySlice_l401_5_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l401_5_4);
  assign _zz_when_ArraySlice_l401_5_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l401_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l401_5_5 = {5'd0, _zz_when_ArraySlice_l401_5_6};
  assign _zz_when_ArraySlice_l401_5_7 = (bReg * 3'b101);
  assign _zz_selectReadFifo_5_15 = 1'b1;
  assign _zz_selectReadFifo_5_14 = {5'd0, _zz_selectReadFifo_5_15};
  assign _zz_when_ArraySlice_l405_5 = (_zz_when_ArraySlice_l405_5_1 % aReg);
  assign _zz_when_ArraySlice_l405_5_1 = (handshakeTimes_5_value + _zz_when_ArraySlice_l405_5_2);
  assign _zz_when_ArraySlice_l405_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l405_5_2 = {12'd0, _zz_when_ArraySlice_l405_5_3};
  assign _zz_when_ArraySlice_l409_5_1 = (selectReadFifo_5 + _zz_when_ArraySlice_l409_5_2);
  assign _zz_when_ArraySlice_l409_5_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l410_5_1 = (_zz_when_ArraySlice_l410_5_2 - _zz_when_ArraySlice_l410_5_3);
  assign _zz_when_ArraySlice_l410_5 = {7'd0, _zz_when_ArraySlice_l410_5_1};
  assign _zz_when_ArraySlice_l410_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l410_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l410_5_3 = {5'd0, _zz_when_ArraySlice_l410_5_4};
  assign _zz__zz_when_ArraySlice_l94_16 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_16 = (_zz_when_ArraySlice_l95_16_1 - _zz_when_ArraySlice_l95_16_4);
  assign _zz_when_ArraySlice_l95_16_1 = (_zz_when_ArraySlice_l95_16_2 + _zz_when_ArraySlice_l95_16_3);
  assign _zz_when_ArraySlice_l95_16_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_16_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_16_4 = {1'd0, _zz_when_ArraySlice_l94_16};
  assign _zz__zz_when_ArraySlice_l412_5 = (_zz__zz_when_ArraySlice_l412_5_1 + _zz__zz_when_ArraySlice_l412_5_2);
  assign _zz__zz_when_ArraySlice_l412_5_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l412_5_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l412_5_3 = {1'd0, _zz_when_ArraySlice_l94_16};
  assign _zz_when_ArraySlice_l99_16_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_16 = _zz_when_ArraySlice_l99_16_1[5:0];
  assign _zz_when_ArraySlice_l412_5_1 = (outSliceNumb_5_value + _zz_when_ArraySlice_l412_5_2);
  assign _zz_when_ArraySlice_l412_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l412_5_2 = {6'd0, _zz_when_ArraySlice_l412_5_3};
  assign _zz_when_ArraySlice_l412_5_4 = (_zz_when_ArraySlice_l412_5 / aReg);
  assign _zz_selectReadFifo_5_16 = (selectReadFifo_5 - _zz_selectReadFifo_5_17);
  assign _zz_selectReadFifo_5_17 = {3'd0, bReg};
  assign _zz_selectReadFifo_5_19 = 1'b1;
  assign _zz_selectReadFifo_5_18 = {5'd0, _zz_selectReadFifo_5_19};
  assign _zz_selectReadFifo_5_20 = (selectReadFifo_5 + _zz_selectReadFifo_5_21);
  assign _zz_selectReadFifo_5_21 = (3'b111 * bReg);
  assign _zz_selectReadFifo_5_23 = 1'b1;
  assign _zz_selectReadFifo_5_22 = {5'd0, _zz_selectReadFifo_5_23};
  assign _zz_when_ArraySlice_l165_136 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_136_1);
  assign _zz_when_ArraySlice_l165_136_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_136_1 = {3'd0, _zz_when_ArraySlice_l165_136_2};
  assign _zz_when_ArraySlice_l166_136 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_136_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_136_3);
  assign _zz_when_ArraySlice_l166_136_1 = {1'd0, _zz_when_ArraySlice_l166_136_2};
  assign _zz_when_ArraySlice_l166_136_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_136_4);
  assign _zz_when_ArraySlice_l166_136_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_136_4 = {3'd0, _zz_when_ArraySlice_l166_136_5};
  assign _zz__zz_when_ArraySlice_l112_136 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_136 = (_zz_when_ArraySlice_l113_136_1 - _zz_when_ArraySlice_l113_136_4);
  assign _zz_when_ArraySlice_l113_136_1 = (_zz_when_ArraySlice_l113_136_2 + _zz_when_ArraySlice_l113_136_3);
  assign _zz_when_ArraySlice_l113_136_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_136_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_136_4 = {1'd0, _zz_when_ArraySlice_l112_136};
  assign _zz__zz_when_ArraySlice_l173_136 = (_zz__zz_when_ArraySlice_l173_136_1 + _zz__zz_when_ArraySlice_l173_136_2);
  assign _zz__zz_when_ArraySlice_l173_136_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_136_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_136_3 = {1'd0, _zz_when_ArraySlice_l112_136};
  assign _zz_when_ArraySlice_l118_136_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_136 = _zz_when_ArraySlice_l118_136_1[5:0];
  assign _zz_when_ArraySlice_l173_136_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_136_2 = (_zz_when_ArraySlice_l173_136_3 + _zz_when_ArraySlice_l173_136_8);
  assign _zz_when_ArraySlice_l173_136_3 = (_zz_when_ArraySlice_l173_136 - _zz_when_ArraySlice_l173_136_4);
  assign _zz_when_ArraySlice_l173_136_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_136_6);
  assign _zz_when_ArraySlice_l173_136_4 = {1'd0, _zz_when_ArraySlice_l173_136_5};
  assign _zz_when_ArraySlice_l173_136_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_136_6 = {3'd0, _zz_when_ArraySlice_l173_136_7};
  assign _zz_when_ArraySlice_l173_136_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_137 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_137_1);
  assign _zz_when_ArraySlice_l165_137_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_137_1 = {2'd0, _zz_when_ArraySlice_l165_137_2};
  assign _zz_when_ArraySlice_l166_137 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_137_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_137_2);
  assign _zz_when_ArraySlice_l166_137_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_137_3);
  assign _zz_when_ArraySlice_l166_137_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_137_3 = {2'd0, _zz_when_ArraySlice_l166_137_4};
  assign _zz__zz_when_ArraySlice_l112_137 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_137 = (_zz_when_ArraySlice_l113_137_1 - _zz_when_ArraySlice_l113_137_4);
  assign _zz_when_ArraySlice_l113_137_1 = (_zz_when_ArraySlice_l113_137_2 + _zz_when_ArraySlice_l113_137_3);
  assign _zz_when_ArraySlice_l113_137_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_137_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_137_4 = {1'd0, _zz_when_ArraySlice_l112_137};
  assign _zz__zz_when_ArraySlice_l173_137 = (_zz__zz_when_ArraySlice_l173_137_1 + _zz__zz_when_ArraySlice_l173_137_2);
  assign _zz__zz_when_ArraySlice_l173_137_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_137_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_137_3 = {1'd0, _zz_when_ArraySlice_l112_137};
  assign _zz_when_ArraySlice_l118_137_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_137 = _zz_when_ArraySlice_l118_137_1[5:0];
  assign _zz_when_ArraySlice_l173_137_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_137_1 = {1'd0, _zz_when_ArraySlice_l173_137_2};
  assign _zz_when_ArraySlice_l173_137_3 = (_zz_when_ArraySlice_l173_137_4 + _zz_when_ArraySlice_l173_137_9);
  assign _zz_when_ArraySlice_l173_137_4 = (_zz_when_ArraySlice_l173_137 - _zz_when_ArraySlice_l173_137_5);
  assign _zz_when_ArraySlice_l173_137_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_137_7);
  assign _zz_when_ArraySlice_l173_137_5 = {1'd0, _zz_when_ArraySlice_l173_137_6};
  assign _zz_when_ArraySlice_l173_137_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_137_7 = {2'd0, _zz_when_ArraySlice_l173_137_8};
  assign _zz_when_ArraySlice_l173_137_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_138 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_138_1);
  assign _zz_when_ArraySlice_l165_138_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_138_1 = {1'd0, _zz_when_ArraySlice_l165_138_2};
  assign _zz_when_ArraySlice_l166_138 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_138_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_138_2);
  assign _zz_when_ArraySlice_l166_138_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_138_3);
  assign _zz_when_ArraySlice_l166_138_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_138_3 = {1'd0, _zz_when_ArraySlice_l166_138_4};
  assign _zz__zz_when_ArraySlice_l112_138 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_138 = (_zz_when_ArraySlice_l113_138_1 - _zz_when_ArraySlice_l113_138_4);
  assign _zz_when_ArraySlice_l113_138_1 = (_zz_when_ArraySlice_l113_138_2 + _zz_when_ArraySlice_l113_138_3);
  assign _zz_when_ArraySlice_l113_138_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_138_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_138_4 = {1'd0, _zz_when_ArraySlice_l112_138};
  assign _zz__zz_when_ArraySlice_l173_138 = (_zz__zz_when_ArraySlice_l173_138_1 + _zz__zz_when_ArraySlice_l173_138_2);
  assign _zz__zz_when_ArraySlice_l173_138_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_138_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_138_3 = {1'd0, _zz_when_ArraySlice_l112_138};
  assign _zz_when_ArraySlice_l118_138_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_138 = _zz_when_ArraySlice_l118_138_1[5:0];
  assign _zz_when_ArraySlice_l173_138_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_138_1 = {1'd0, _zz_when_ArraySlice_l173_138_2};
  assign _zz_when_ArraySlice_l173_138_3 = (_zz_when_ArraySlice_l173_138_4 + _zz_when_ArraySlice_l173_138_9);
  assign _zz_when_ArraySlice_l173_138_4 = (_zz_when_ArraySlice_l173_138 - _zz_when_ArraySlice_l173_138_5);
  assign _zz_when_ArraySlice_l173_138_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_138_7);
  assign _zz_when_ArraySlice_l173_138_5 = {1'd0, _zz_when_ArraySlice_l173_138_6};
  assign _zz_when_ArraySlice_l173_138_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_138_7 = {1'd0, _zz_when_ArraySlice_l173_138_8};
  assign _zz_when_ArraySlice_l173_138_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_139 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_139_1);
  assign _zz_when_ArraySlice_l165_139_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_139_1 = {1'd0, _zz_when_ArraySlice_l165_139_2};
  assign _zz_when_ArraySlice_l166_139 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_139_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_139_2);
  assign _zz_when_ArraySlice_l166_139_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_139_3);
  assign _zz_when_ArraySlice_l166_139_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_139_3 = {1'd0, _zz_when_ArraySlice_l166_139_4};
  assign _zz__zz_when_ArraySlice_l112_139 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_139 = (_zz_when_ArraySlice_l113_139_1 - _zz_when_ArraySlice_l113_139_4);
  assign _zz_when_ArraySlice_l113_139_1 = (_zz_when_ArraySlice_l113_139_2 + _zz_when_ArraySlice_l113_139_3);
  assign _zz_when_ArraySlice_l113_139_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_139_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_139_4 = {1'd0, _zz_when_ArraySlice_l112_139};
  assign _zz__zz_when_ArraySlice_l173_139 = (_zz__zz_when_ArraySlice_l173_139_1 + _zz__zz_when_ArraySlice_l173_139_2);
  assign _zz__zz_when_ArraySlice_l173_139_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_139_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_139_3 = {1'd0, _zz_when_ArraySlice_l112_139};
  assign _zz_when_ArraySlice_l118_139_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_139 = _zz_when_ArraySlice_l118_139_1[5:0];
  assign _zz_when_ArraySlice_l173_139_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_139_1 = {1'd0, _zz_when_ArraySlice_l173_139_2};
  assign _zz_when_ArraySlice_l173_139_3 = (_zz_when_ArraySlice_l173_139_4 + _zz_when_ArraySlice_l173_139_9);
  assign _zz_when_ArraySlice_l173_139_4 = (_zz_when_ArraySlice_l173_139 - _zz_when_ArraySlice_l173_139_5);
  assign _zz_when_ArraySlice_l173_139_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_139_7);
  assign _zz_when_ArraySlice_l173_139_5 = {1'd0, _zz_when_ArraySlice_l173_139_6};
  assign _zz_when_ArraySlice_l173_139_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_139_7 = {1'd0, _zz_when_ArraySlice_l173_139_8};
  assign _zz_when_ArraySlice_l173_139_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_140 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_140_1);
  assign _zz_when_ArraySlice_l165_140_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_140 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_140_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_140_2);
  assign _zz_when_ArraySlice_l166_140_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_140_3);
  assign _zz_when_ArraySlice_l166_140_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_140 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_140 = (_zz_when_ArraySlice_l113_140_1 - _zz_when_ArraySlice_l113_140_4);
  assign _zz_when_ArraySlice_l113_140_1 = (_zz_when_ArraySlice_l113_140_2 + _zz_when_ArraySlice_l113_140_3);
  assign _zz_when_ArraySlice_l113_140_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_140_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_140_4 = {1'd0, _zz_when_ArraySlice_l112_140};
  assign _zz__zz_when_ArraySlice_l173_140 = (_zz__zz_when_ArraySlice_l173_140_1 + _zz__zz_when_ArraySlice_l173_140_2);
  assign _zz__zz_when_ArraySlice_l173_140_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_140_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_140_3 = {1'd0, _zz_when_ArraySlice_l112_140};
  assign _zz_when_ArraySlice_l118_140_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_140 = _zz_when_ArraySlice_l118_140_1[5:0];
  assign _zz_when_ArraySlice_l173_140_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_140_1 = {1'd0, _zz_when_ArraySlice_l173_140_2};
  assign _zz_when_ArraySlice_l173_140_3 = (_zz_when_ArraySlice_l173_140_4 + _zz_when_ArraySlice_l173_140_8);
  assign _zz_when_ArraySlice_l173_140_4 = (_zz_when_ArraySlice_l173_140 - _zz_when_ArraySlice_l173_140_5);
  assign _zz_when_ArraySlice_l173_140_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_140_7);
  assign _zz_when_ArraySlice_l173_140_5 = {1'd0, _zz_when_ArraySlice_l173_140_6};
  assign _zz_when_ArraySlice_l173_140_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_140_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_141 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_141_1);
  assign _zz_when_ArraySlice_l165_141_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_141_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_141 = {1'd0, _zz_when_ArraySlice_l166_141_1};
  assign _zz_when_ArraySlice_l166_141_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_141_3);
  assign _zz_when_ArraySlice_l166_141_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_141_4);
  assign _zz_when_ArraySlice_l166_141_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_141 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_141 = (_zz_when_ArraySlice_l113_141_1 - _zz_when_ArraySlice_l113_141_4);
  assign _zz_when_ArraySlice_l113_141_1 = (_zz_when_ArraySlice_l113_141_2 + _zz_when_ArraySlice_l113_141_3);
  assign _zz_when_ArraySlice_l113_141_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_141_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_141_4 = {1'd0, _zz_when_ArraySlice_l112_141};
  assign _zz__zz_when_ArraySlice_l173_141 = (_zz__zz_when_ArraySlice_l173_141_1 + _zz__zz_when_ArraySlice_l173_141_2);
  assign _zz__zz_when_ArraySlice_l173_141_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_141_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_141_3 = {1'd0, _zz_when_ArraySlice_l112_141};
  assign _zz_when_ArraySlice_l118_141_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_141 = _zz_when_ArraySlice_l118_141_1[5:0];
  assign _zz_when_ArraySlice_l173_141_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_141_1 = {2'd0, _zz_when_ArraySlice_l173_141_2};
  assign _zz_when_ArraySlice_l173_141_3 = (_zz_when_ArraySlice_l173_141_4 + _zz_when_ArraySlice_l173_141_8);
  assign _zz_when_ArraySlice_l173_141_4 = (_zz_when_ArraySlice_l173_141 - _zz_when_ArraySlice_l173_141_5);
  assign _zz_when_ArraySlice_l173_141_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_141_7);
  assign _zz_when_ArraySlice_l173_141_5 = {1'd0, _zz_when_ArraySlice_l173_141_6};
  assign _zz_when_ArraySlice_l173_141_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_141_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_142 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_142_1);
  assign _zz_when_ArraySlice_l165_142_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_142_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_142 = {1'd0, _zz_when_ArraySlice_l166_142_1};
  assign _zz_when_ArraySlice_l166_142_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_142_3);
  assign _zz_when_ArraySlice_l166_142_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_142_4);
  assign _zz_when_ArraySlice_l166_142_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_142 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_142 = (_zz_when_ArraySlice_l113_142_1 - _zz_when_ArraySlice_l113_142_4);
  assign _zz_when_ArraySlice_l113_142_1 = (_zz_when_ArraySlice_l113_142_2 + _zz_when_ArraySlice_l113_142_3);
  assign _zz_when_ArraySlice_l113_142_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_142_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_142_4 = {1'd0, _zz_when_ArraySlice_l112_142};
  assign _zz__zz_when_ArraySlice_l173_142 = (_zz__zz_when_ArraySlice_l173_142_1 + _zz__zz_when_ArraySlice_l173_142_2);
  assign _zz__zz_when_ArraySlice_l173_142_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_142_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_142_3 = {1'd0, _zz_when_ArraySlice_l112_142};
  assign _zz_when_ArraySlice_l118_142_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_142 = _zz_when_ArraySlice_l118_142_1[5:0];
  assign _zz_when_ArraySlice_l173_142_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_142_1 = {2'd0, _zz_when_ArraySlice_l173_142_2};
  assign _zz_when_ArraySlice_l173_142_3 = (_zz_when_ArraySlice_l173_142_4 + _zz_when_ArraySlice_l173_142_8);
  assign _zz_when_ArraySlice_l173_142_4 = (_zz_when_ArraySlice_l173_142 - _zz_when_ArraySlice_l173_142_5);
  assign _zz_when_ArraySlice_l173_142_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_142_7);
  assign _zz_when_ArraySlice_l173_142_5 = {1'd0, _zz_when_ArraySlice_l173_142_6};
  assign _zz_when_ArraySlice_l173_142_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_142_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_143 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_143_1);
  assign _zz_when_ArraySlice_l165_143_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_143_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_143 = {2'd0, _zz_when_ArraySlice_l166_143_1};
  assign _zz_when_ArraySlice_l166_143_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_143_3);
  assign _zz_when_ArraySlice_l166_143_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_143_4);
  assign _zz_when_ArraySlice_l166_143_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_143 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_143 = (_zz_when_ArraySlice_l113_143_1 - _zz_when_ArraySlice_l113_143_4);
  assign _zz_when_ArraySlice_l113_143_1 = (_zz_when_ArraySlice_l113_143_2 + _zz_when_ArraySlice_l113_143_3);
  assign _zz_when_ArraySlice_l113_143_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_143_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_143_4 = {1'd0, _zz_when_ArraySlice_l112_143};
  assign _zz__zz_when_ArraySlice_l173_143 = (_zz__zz_when_ArraySlice_l173_143_1 + _zz__zz_when_ArraySlice_l173_143_2);
  assign _zz__zz_when_ArraySlice_l173_143_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_143_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_143_3 = {1'd0, _zz_when_ArraySlice_l112_143};
  assign _zz_when_ArraySlice_l118_143_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_143 = _zz_when_ArraySlice_l118_143_1[5:0];
  assign _zz_when_ArraySlice_l173_143_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_143_1 = {3'd0, _zz_when_ArraySlice_l173_143_2};
  assign _zz_when_ArraySlice_l173_143_3 = (_zz_when_ArraySlice_l173_143_4 + _zz_when_ArraySlice_l173_143_8);
  assign _zz_when_ArraySlice_l173_143_4 = (_zz_when_ArraySlice_l173_143 - _zz_when_ArraySlice_l173_143_5);
  assign _zz_when_ArraySlice_l173_143_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_143_7);
  assign _zz_when_ArraySlice_l173_143_5 = {1'd0, _zz_when_ArraySlice_l173_143_6};
  assign _zz_when_ArraySlice_l173_143_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_143_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l421_5_1 = (_zz_when_ArraySlice_l421_5_2 + _zz_when_ArraySlice_l421_5_7);
  assign _zz_when_ArraySlice_l421_5_2 = (_zz_when_ArraySlice_l421_5_3 + _zz_when_ArraySlice_l421_5_5);
  assign _zz_when_ArraySlice_l421_5_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l421_5_4);
  assign _zz_when_ArraySlice_l421_5_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l421_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l421_5_5 = {5'd0, _zz_when_ArraySlice_l421_5_6};
  assign _zz_when_ArraySlice_l421_5_7 = (bReg * 3'b101);
  assign _zz_selectReadFifo_5_25 = 1'b1;
  assign _zz_selectReadFifo_5_24 = {5'd0, _zz_selectReadFifo_5_25};
  assign _zz_when_ArraySlice_l425_5 = (_zz_when_ArraySlice_l425_5_1 % aReg);
  assign _zz_when_ArraySlice_l425_5_1 = (handshakeTimes_5_value + _zz_when_ArraySlice_l425_5_2);
  assign _zz_when_ArraySlice_l425_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l425_5_2 = {12'd0, _zz_when_ArraySlice_l425_5_3};
  assign _zz_when_ArraySlice_l436_5_1 = (_zz_when_ArraySlice_l436_5_2 - _zz_when_ArraySlice_l436_5_3);
  assign _zz_when_ArraySlice_l436_5 = {7'd0, _zz_when_ArraySlice_l436_5_1};
  assign _zz_when_ArraySlice_l436_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l436_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l436_5_3 = {5'd0, _zz_when_ArraySlice_l436_5_4};
  assign _zz__zz_when_ArraySlice_l94_17 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_17 = (_zz_when_ArraySlice_l95_17_1 - _zz_when_ArraySlice_l95_17_4);
  assign _zz_when_ArraySlice_l95_17_1 = (_zz_when_ArraySlice_l95_17_2 + _zz_when_ArraySlice_l95_17_3);
  assign _zz_when_ArraySlice_l95_17_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_17_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_17_4 = {1'd0, _zz_when_ArraySlice_l94_17};
  assign _zz__zz_when_ArraySlice_l437_5 = (_zz__zz_when_ArraySlice_l437_5_1 + _zz__zz_when_ArraySlice_l437_5_2);
  assign _zz__zz_when_ArraySlice_l437_5_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l437_5_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l437_5_3 = {1'd0, _zz_when_ArraySlice_l94_17};
  assign _zz_when_ArraySlice_l99_17_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_17 = _zz_when_ArraySlice_l99_17_1[5:0];
  assign _zz_when_ArraySlice_l437_5_1 = (outSliceNumb_5_value + _zz_when_ArraySlice_l437_5_2);
  assign _zz_when_ArraySlice_l437_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l437_5_2 = {6'd0, _zz_when_ArraySlice_l437_5_3};
  assign _zz_when_ArraySlice_l437_5_4 = (_zz_when_ArraySlice_l437_5 / aReg);
  assign _zz_selectReadFifo_5_26 = (selectReadFifo_5 - _zz_selectReadFifo_5_27);
  assign _zz_selectReadFifo_5_27 = {3'd0, bReg};
  assign _zz_selectReadFifo_5_29 = 1'b1;
  assign _zz_selectReadFifo_5_28 = {5'd0, _zz_selectReadFifo_5_29};
  assign _zz_when_ArraySlice_l165_144 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_144_1);
  assign _zz_when_ArraySlice_l165_144_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_144_1 = {3'd0, _zz_when_ArraySlice_l165_144_2};
  assign _zz_when_ArraySlice_l166_144 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_144_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_144_3);
  assign _zz_when_ArraySlice_l166_144_1 = {1'd0, _zz_when_ArraySlice_l166_144_2};
  assign _zz_when_ArraySlice_l166_144_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_144_4);
  assign _zz_when_ArraySlice_l166_144_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_144_4 = {3'd0, _zz_when_ArraySlice_l166_144_5};
  assign _zz__zz_when_ArraySlice_l112_144 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_144 = (_zz_when_ArraySlice_l113_144_1 - _zz_when_ArraySlice_l113_144_4);
  assign _zz_when_ArraySlice_l113_144_1 = (_zz_when_ArraySlice_l113_144_2 + _zz_when_ArraySlice_l113_144_3);
  assign _zz_when_ArraySlice_l113_144_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_144_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_144_4 = {1'd0, _zz_when_ArraySlice_l112_144};
  assign _zz__zz_when_ArraySlice_l173_144 = (_zz__zz_when_ArraySlice_l173_144_1 + _zz__zz_when_ArraySlice_l173_144_2);
  assign _zz__zz_when_ArraySlice_l173_144_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_144_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_144_3 = {1'd0, _zz_when_ArraySlice_l112_144};
  assign _zz_when_ArraySlice_l118_144_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_144 = _zz_when_ArraySlice_l118_144_1[5:0];
  assign _zz_when_ArraySlice_l173_144_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_144_2 = (_zz_when_ArraySlice_l173_144_3 + _zz_when_ArraySlice_l173_144_8);
  assign _zz_when_ArraySlice_l173_144_3 = (_zz_when_ArraySlice_l173_144 - _zz_when_ArraySlice_l173_144_4);
  assign _zz_when_ArraySlice_l173_144_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_144_6);
  assign _zz_when_ArraySlice_l173_144_4 = {1'd0, _zz_when_ArraySlice_l173_144_5};
  assign _zz_when_ArraySlice_l173_144_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_144_6 = {3'd0, _zz_when_ArraySlice_l173_144_7};
  assign _zz_when_ArraySlice_l173_144_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_145 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_145_1);
  assign _zz_when_ArraySlice_l165_145_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_145_1 = {2'd0, _zz_when_ArraySlice_l165_145_2};
  assign _zz_when_ArraySlice_l166_145 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_145_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_145_2);
  assign _zz_when_ArraySlice_l166_145_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_145_3);
  assign _zz_when_ArraySlice_l166_145_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_145_3 = {2'd0, _zz_when_ArraySlice_l166_145_4};
  assign _zz__zz_when_ArraySlice_l112_145 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_145 = (_zz_when_ArraySlice_l113_145_1 - _zz_when_ArraySlice_l113_145_4);
  assign _zz_when_ArraySlice_l113_145_1 = (_zz_when_ArraySlice_l113_145_2 + _zz_when_ArraySlice_l113_145_3);
  assign _zz_when_ArraySlice_l113_145_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_145_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_145_4 = {1'd0, _zz_when_ArraySlice_l112_145};
  assign _zz__zz_when_ArraySlice_l173_145 = (_zz__zz_when_ArraySlice_l173_145_1 + _zz__zz_when_ArraySlice_l173_145_2);
  assign _zz__zz_when_ArraySlice_l173_145_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_145_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_145_3 = {1'd0, _zz_when_ArraySlice_l112_145};
  assign _zz_when_ArraySlice_l118_145_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_145 = _zz_when_ArraySlice_l118_145_1[5:0];
  assign _zz_when_ArraySlice_l173_145_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_145_1 = {1'd0, _zz_when_ArraySlice_l173_145_2};
  assign _zz_when_ArraySlice_l173_145_3 = (_zz_when_ArraySlice_l173_145_4 + _zz_when_ArraySlice_l173_145_9);
  assign _zz_when_ArraySlice_l173_145_4 = (_zz_when_ArraySlice_l173_145 - _zz_when_ArraySlice_l173_145_5);
  assign _zz_when_ArraySlice_l173_145_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_145_7);
  assign _zz_when_ArraySlice_l173_145_5 = {1'd0, _zz_when_ArraySlice_l173_145_6};
  assign _zz_when_ArraySlice_l173_145_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_145_7 = {2'd0, _zz_when_ArraySlice_l173_145_8};
  assign _zz_when_ArraySlice_l173_145_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_146 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_146_1);
  assign _zz_when_ArraySlice_l165_146_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_146_1 = {1'd0, _zz_when_ArraySlice_l165_146_2};
  assign _zz_when_ArraySlice_l166_146 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_146_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_146_2);
  assign _zz_when_ArraySlice_l166_146_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_146_3);
  assign _zz_when_ArraySlice_l166_146_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_146_3 = {1'd0, _zz_when_ArraySlice_l166_146_4};
  assign _zz__zz_when_ArraySlice_l112_146 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_146 = (_zz_when_ArraySlice_l113_146_1 - _zz_when_ArraySlice_l113_146_4);
  assign _zz_when_ArraySlice_l113_146_1 = (_zz_when_ArraySlice_l113_146_2 + _zz_when_ArraySlice_l113_146_3);
  assign _zz_when_ArraySlice_l113_146_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_146_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_146_4 = {1'd0, _zz_when_ArraySlice_l112_146};
  assign _zz__zz_when_ArraySlice_l173_146 = (_zz__zz_when_ArraySlice_l173_146_1 + _zz__zz_when_ArraySlice_l173_146_2);
  assign _zz__zz_when_ArraySlice_l173_146_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_146_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_146_3 = {1'd0, _zz_when_ArraySlice_l112_146};
  assign _zz_when_ArraySlice_l118_146_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_146 = _zz_when_ArraySlice_l118_146_1[5:0];
  assign _zz_when_ArraySlice_l173_146_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_146_1 = {1'd0, _zz_when_ArraySlice_l173_146_2};
  assign _zz_when_ArraySlice_l173_146_3 = (_zz_when_ArraySlice_l173_146_4 + _zz_when_ArraySlice_l173_146_9);
  assign _zz_when_ArraySlice_l173_146_4 = (_zz_when_ArraySlice_l173_146 - _zz_when_ArraySlice_l173_146_5);
  assign _zz_when_ArraySlice_l173_146_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_146_7);
  assign _zz_when_ArraySlice_l173_146_5 = {1'd0, _zz_when_ArraySlice_l173_146_6};
  assign _zz_when_ArraySlice_l173_146_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_146_7 = {1'd0, _zz_when_ArraySlice_l173_146_8};
  assign _zz_when_ArraySlice_l173_146_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_147 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_147_1);
  assign _zz_when_ArraySlice_l165_147_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_147_1 = {1'd0, _zz_when_ArraySlice_l165_147_2};
  assign _zz_when_ArraySlice_l166_147 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_147_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_147_2);
  assign _zz_when_ArraySlice_l166_147_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_147_3);
  assign _zz_when_ArraySlice_l166_147_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_147_3 = {1'd0, _zz_when_ArraySlice_l166_147_4};
  assign _zz__zz_when_ArraySlice_l112_147 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_147 = (_zz_when_ArraySlice_l113_147_1 - _zz_when_ArraySlice_l113_147_4);
  assign _zz_when_ArraySlice_l113_147_1 = (_zz_when_ArraySlice_l113_147_2 + _zz_when_ArraySlice_l113_147_3);
  assign _zz_when_ArraySlice_l113_147_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_147_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_147_4 = {1'd0, _zz_when_ArraySlice_l112_147};
  assign _zz__zz_when_ArraySlice_l173_147 = (_zz__zz_when_ArraySlice_l173_147_1 + _zz__zz_when_ArraySlice_l173_147_2);
  assign _zz__zz_when_ArraySlice_l173_147_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_147_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_147_3 = {1'd0, _zz_when_ArraySlice_l112_147};
  assign _zz_when_ArraySlice_l118_147_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_147 = _zz_when_ArraySlice_l118_147_1[5:0];
  assign _zz_when_ArraySlice_l173_147_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_147_1 = {1'd0, _zz_when_ArraySlice_l173_147_2};
  assign _zz_when_ArraySlice_l173_147_3 = (_zz_when_ArraySlice_l173_147_4 + _zz_when_ArraySlice_l173_147_9);
  assign _zz_when_ArraySlice_l173_147_4 = (_zz_when_ArraySlice_l173_147 - _zz_when_ArraySlice_l173_147_5);
  assign _zz_when_ArraySlice_l173_147_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_147_7);
  assign _zz_when_ArraySlice_l173_147_5 = {1'd0, _zz_when_ArraySlice_l173_147_6};
  assign _zz_when_ArraySlice_l173_147_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_147_7 = {1'd0, _zz_when_ArraySlice_l173_147_8};
  assign _zz_when_ArraySlice_l173_147_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_148 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_148_1);
  assign _zz_when_ArraySlice_l165_148_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_148 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_148_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_148_2);
  assign _zz_when_ArraySlice_l166_148_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_148_3);
  assign _zz_when_ArraySlice_l166_148_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_148 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_148 = (_zz_when_ArraySlice_l113_148_1 - _zz_when_ArraySlice_l113_148_4);
  assign _zz_when_ArraySlice_l113_148_1 = (_zz_when_ArraySlice_l113_148_2 + _zz_when_ArraySlice_l113_148_3);
  assign _zz_when_ArraySlice_l113_148_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_148_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_148_4 = {1'd0, _zz_when_ArraySlice_l112_148};
  assign _zz__zz_when_ArraySlice_l173_148 = (_zz__zz_when_ArraySlice_l173_148_1 + _zz__zz_when_ArraySlice_l173_148_2);
  assign _zz__zz_when_ArraySlice_l173_148_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_148_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_148_3 = {1'd0, _zz_when_ArraySlice_l112_148};
  assign _zz_when_ArraySlice_l118_148_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_148 = _zz_when_ArraySlice_l118_148_1[5:0];
  assign _zz_when_ArraySlice_l173_148_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_148_1 = {1'd0, _zz_when_ArraySlice_l173_148_2};
  assign _zz_when_ArraySlice_l173_148_3 = (_zz_when_ArraySlice_l173_148_4 + _zz_when_ArraySlice_l173_148_8);
  assign _zz_when_ArraySlice_l173_148_4 = (_zz_when_ArraySlice_l173_148 - _zz_when_ArraySlice_l173_148_5);
  assign _zz_when_ArraySlice_l173_148_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_148_7);
  assign _zz_when_ArraySlice_l173_148_5 = {1'd0, _zz_when_ArraySlice_l173_148_6};
  assign _zz_when_ArraySlice_l173_148_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_148_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_149 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_149_1);
  assign _zz_when_ArraySlice_l165_149_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_149_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_149 = {1'd0, _zz_when_ArraySlice_l166_149_1};
  assign _zz_when_ArraySlice_l166_149_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_149_3);
  assign _zz_when_ArraySlice_l166_149_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_149_4);
  assign _zz_when_ArraySlice_l166_149_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_149 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_149 = (_zz_when_ArraySlice_l113_149_1 - _zz_when_ArraySlice_l113_149_4);
  assign _zz_when_ArraySlice_l113_149_1 = (_zz_when_ArraySlice_l113_149_2 + _zz_when_ArraySlice_l113_149_3);
  assign _zz_when_ArraySlice_l113_149_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_149_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_149_4 = {1'd0, _zz_when_ArraySlice_l112_149};
  assign _zz__zz_when_ArraySlice_l173_149 = (_zz__zz_when_ArraySlice_l173_149_1 + _zz__zz_when_ArraySlice_l173_149_2);
  assign _zz__zz_when_ArraySlice_l173_149_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_149_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_149_3 = {1'd0, _zz_when_ArraySlice_l112_149};
  assign _zz_when_ArraySlice_l118_149_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_149 = _zz_when_ArraySlice_l118_149_1[5:0];
  assign _zz_when_ArraySlice_l173_149_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_149_1 = {2'd0, _zz_when_ArraySlice_l173_149_2};
  assign _zz_when_ArraySlice_l173_149_3 = (_zz_when_ArraySlice_l173_149_4 + _zz_when_ArraySlice_l173_149_8);
  assign _zz_when_ArraySlice_l173_149_4 = (_zz_when_ArraySlice_l173_149 - _zz_when_ArraySlice_l173_149_5);
  assign _zz_when_ArraySlice_l173_149_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_149_7);
  assign _zz_when_ArraySlice_l173_149_5 = {1'd0, _zz_when_ArraySlice_l173_149_6};
  assign _zz_when_ArraySlice_l173_149_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_149_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_150 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_150_1);
  assign _zz_when_ArraySlice_l165_150_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_150_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_150 = {1'd0, _zz_when_ArraySlice_l166_150_1};
  assign _zz_when_ArraySlice_l166_150_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_150_3);
  assign _zz_when_ArraySlice_l166_150_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_150_4);
  assign _zz_when_ArraySlice_l166_150_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_150 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_150 = (_zz_when_ArraySlice_l113_150_1 - _zz_when_ArraySlice_l113_150_4);
  assign _zz_when_ArraySlice_l113_150_1 = (_zz_when_ArraySlice_l113_150_2 + _zz_when_ArraySlice_l113_150_3);
  assign _zz_when_ArraySlice_l113_150_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_150_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_150_4 = {1'd0, _zz_when_ArraySlice_l112_150};
  assign _zz__zz_when_ArraySlice_l173_150 = (_zz__zz_when_ArraySlice_l173_150_1 + _zz__zz_when_ArraySlice_l173_150_2);
  assign _zz__zz_when_ArraySlice_l173_150_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_150_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_150_3 = {1'd0, _zz_when_ArraySlice_l112_150};
  assign _zz_when_ArraySlice_l118_150_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_150 = _zz_when_ArraySlice_l118_150_1[5:0];
  assign _zz_when_ArraySlice_l173_150_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_150_1 = {2'd0, _zz_when_ArraySlice_l173_150_2};
  assign _zz_when_ArraySlice_l173_150_3 = (_zz_when_ArraySlice_l173_150_4 + _zz_when_ArraySlice_l173_150_8);
  assign _zz_when_ArraySlice_l173_150_4 = (_zz_when_ArraySlice_l173_150 - _zz_when_ArraySlice_l173_150_5);
  assign _zz_when_ArraySlice_l173_150_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_150_7);
  assign _zz_when_ArraySlice_l173_150_5 = {1'd0, _zz_when_ArraySlice_l173_150_6};
  assign _zz_when_ArraySlice_l173_150_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_150_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_151 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_151_1);
  assign _zz_when_ArraySlice_l165_151_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_151_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_151 = {2'd0, _zz_when_ArraySlice_l166_151_1};
  assign _zz_when_ArraySlice_l166_151_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_151_3);
  assign _zz_when_ArraySlice_l166_151_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_151_4);
  assign _zz_when_ArraySlice_l166_151_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_151 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_151 = (_zz_when_ArraySlice_l113_151_1 - _zz_when_ArraySlice_l113_151_4);
  assign _zz_when_ArraySlice_l113_151_1 = (_zz_when_ArraySlice_l113_151_2 + _zz_when_ArraySlice_l113_151_3);
  assign _zz_when_ArraySlice_l113_151_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_151_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_151_4 = {1'd0, _zz_when_ArraySlice_l112_151};
  assign _zz__zz_when_ArraySlice_l173_151 = (_zz__zz_when_ArraySlice_l173_151_1 + _zz__zz_when_ArraySlice_l173_151_2);
  assign _zz__zz_when_ArraySlice_l173_151_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_151_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_151_3 = {1'd0, _zz_when_ArraySlice_l112_151};
  assign _zz_when_ArraySlice_l118_151_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_151 = _zz_when_ArraySlice_l118_151_1[5:0];
  assign _zz_when_ArraySlice_l173_151_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_151_1 = {3'd0, _zz_when_ArraySlice_l173_151_2};
  assign _zz_when_ArraySlice_l173_151_3 = (_zz_when_ArraySlice_l173_151_4 + _zz_when_ArraySlice_l173_151_8);
  assign _zz_when_ArraySlice_l173_151_4 = (_zz_when_ArraySlice_l173_151 - _zz_when_ArraySlice_l173_151_5);
  assign _zz_when_ArraySlice_l173_151_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_151_7);
  assign _zz_when_ArraySlice_l173_151_5 = {1'd0, _zz_when_ArraySlice_l173_151_6};
  assign _zz_when_ArraySlice_l173_151_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_151_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_5_31 = 1'b1;
  assign _zz_selectReadFifo_5_30 = {5'd0, _zz_selectReadFifo_5_31};
  assign _zz_when_ArraySlice_l448_5 = (_zz_when_ArraySlice_l448_5_1 % aReg);
  assign _zz_when_ArraySlice_l448_5_1 = (handshakeTimes_5_value + _zz_when_ArraySlice_l448_5_2);
  assign _zz_when_ArraySlice_l448_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l448_5_2 = {12'd0, _zz_when_ArraySlice_l448_5_3};
  assign _zz_when_ArraySlice_l434_5 = (selectReadFifo_5 + _zz_when_ArraySlice_l434_5_1);
  assign _zz_when_ArraySlice_l434_5_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l455_5_1 = (_zz_when_ArraySlice_l455_5_2 - _zz_when_ArraySlice_l455_5_3);
  assign _zz_when_ArraySlice_l455_5 = {7'd0, _zz_when_ArraySlice_l455_5_1};
  assign _zz_when_ArraySlice_l455_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l455_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l455_5_3 = {5'd0, _zz_when_ArraySlice_l455_5_4};
  assign _zz_when_ArraySlice_l373_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l373_6_1);
  assign _zz_when_ArraySlice_l373_6_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l374_6_1 = (selectReadFifo_6 + _zz_when_ArraySlice_l374_6_2);
  assign _zz_when_ArraySlice_l374_6_2 = (bReg * 3'b110);
  assign _zz__zz_outputStreamArrayData_6_valid = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l380_6_1 = 1'b1;
  assign _zz_when_ArraySlice_l380_6 = {6'd0, _zz_when_ArraySlice_l380_6_1};
  assign _zz_when_ArraySlice_l380_6_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l380_6_4);
  assign _zz_when_ArraySlice_l380_6_4 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l381_6_1 = (_zz_when_ArraySlice_l381_6_2 - _zz_when_ArraySlice_l381_6_3);
  assign _zz_when_ArraySlice_l381_6 = {7'd0, _zz_when_ArraySlice_l381_6_1};
  assign _zz_when_ArraySlice_l381_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l381_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l381_6_3 = {5'd0, _zz_when_ArraySlice_l381_6_4};
  assign _zz_selectReadFifo_6 = (selectReadFifo_6 - _zz_selectReadFifo_6_1);
  assign _zz_selectReadFifo_6_1 = {3'd0, bReg};
  assign _zz_selectReadFifo_6_3 = 1'b1;
  assign _zz_selectReadFifo_6_2 = {5'd0, _zz_selectReadFifo_6_3};
  assign _zz_selectReadFifo_6_5 = 1'b1;
  assign _zz_selectReadFifo_6_4 = {5'd0, _zz_selectReadFifo_6_5};
  assign _zz_when_ArraySlice_l384_6 = (_zz_when_ArraySlice_l384_6_1 % aReg);
  assign _zz_when_ArraySlice_l384_6_1 = (handshakeTimes_6_value + _zz_when_ArraySlice_l384_6_2);
  assign _zz_when_ArraySlice_l384_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l384_6_2 = {12'd0, _zz_when_ArraySlice_l384_6_3};
  assign _zz_when_ArraySlice_l389_6_1 = (selectReadFifo_6 + _zz_when_ArraySlice_l389_6_2);
  assign _zz_when_ArraySlice_l389_6_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l389_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l389_6_3 = {6'd0, _zz_when_ArraySlice_l389_6_4};
  assign _zz_when_ArraySlice_l390_6_1 = (_zz_when_ArraySlice_l390_6_2 - _zz_when_ArraySlice_l390_6_3);
  assign _zz_when_ArraySlice_l390_6 = {7'd0, _zz_when_ArraySlice_l390_6_1};
  assign _zz_when_ArraySlice_l390_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l390_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l390_6_3 = {5'd0, _zz_when_ArraySlice_l390_6_4};
  assign _zz__zz_when_ArraySlice_l94_18 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_18 = (_zz_when_ArraySlice_l95_18_1 - _zz_when_ArraySlice_l95_18_4);
  assign _zz_when_ArraySlice_l95_18_1 = (_zz_when_ArraySlice_l95_18_2 + _zz_when_ArraySlice_l95_18_3);
  assign _zz_when_ArraySlice_l95_18_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_18_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_18_4 = {1'd0, _zz_when_ArraySlice_l94_18};
  assign _zz__zz_when_ArraySlice_l392_6 = (_zz__zz_when_ArraySlice_l392_6_1 + _zz__zz_when_ArraySlice_l392_6_2);
  assign _zz__zz_when_ArraySlice_l392_6_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l392_6_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l392_6_3 = {1'd0, _zz_when_ArraySlice_l94_18};
  assign _zz_when_ArraySlice_l99_18_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_18 = _zz_when_ArraySlice_l99_18_1[5:0];
  assign _zz_when_ArraySlice_l392_6_1 = (outSliceNumb_6_value + _zz_when_ArraySlice_l392_6_2);
  assign _zz_when_ArraySlice_l392_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l392_6_2 = {6'd0, _zz_when_ArraySlice_l392_6_3};
  assign _zz_when_ArraySlice_l392_6_4 = (_zz_when_ArraySlice_l392_6 / aReg);
  assign _zz_selectReadFifo_6_6 = (selectReadFifo_6 - _zz_selectReadFifo_6_7);
  assign _zz_selectReadFifo_6_7 = {3'd0, bReg};
  assign _zz_selectReadFifo_6_9 = 1'b1;
  assign _zz_selectReadFifo_6_8 = {5'd0, _zz_selectReadFifo_6_9};
  assign _zz_selectReadFifo_6_10 = (selectReadFifo_6 + _zz_selectReadFifo_6_11);
  assign _zz_selectReadFifo_6_11 = (3'b111 * bReg);
  assign _zz_selectReadFifo_6_13 = 1'b1;
  assign _zz_selectReadFifo_6_12 = {5'd0, _zz_selectReadFifo_6_13};
  assign _zz_when_ArraySlice_l165_152 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_152_1);
  assign _zz_when_ArraySlice_l165_152_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_152_1 = {3'd0, _zz_when_ArraySlice_l165_152_2};
  assign _zz_when_ArraySlice_l166_152 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_152_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_152_3);
  assign _zz_when_ArraySlice_l166_152_1 = {1'd0, _zz_when_ArraySlice_l166_152_2};
  assign _zz_when_ArraySlice_l166_152_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_152_4);
  assign _zz_when_ArraySlice_l166_152_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_152_4 = {3'd0, _zz_when_ArraySlice_l166_152_5};
  assign _zz__zz_when_ArraySlice_l112_152 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_152 = (_zz_when_ArraySlice_l113_152_1 - _zz_when_ArraySlice_l113_152_4);
  assign _zz_when_ArraySlice_l113_152_1 = (_zz_when_ArraySlice_l113_152_2 + _zz_when_ArraySlice_l113_152_3);
  assign _zz_when_ArraySlice_l113_152_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_152_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_152_4 = {1'd0, _zz_when_ArraySlice_l112_152};
  assign _zz__zz_when_ArraySlice_l173_152 = (_zz__zz_when_ArraySlice_l173_152_1 + _zz__zz_when_ArraySlice_l173_152_2);
  assign _zz__zz_when_ArraySlice_l173_152_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_152_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_152_3 = {1'd0, _zz_when_ArraySlice_l112_152};
  assign _zz_when_ArraySlice_l118_152_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_152 = _zz_when_ArraySlice_l118_152_1[5:0];
  assign _zz_when_ArraySlice_l173_152_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_152_2 = (_zz_when_ArraySlice_l173_152_3 + _zz_when_ArraySlice_l173_152_8);
  assign _zz_when_ArraySlice_l173_152_3 = (_zz_when_ArraySlice_l173_152 - _zz_when_ArraySlice_l173_152_4);
  assign _zz_when_ArraySlice_l173_152_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_152_6);
  assign _zz_when_ArraySlice_l173_152_4 = {1'd0, _zz_when_ArraySlice_l173_152_5};
  assign _zz_when_ArraySlice_l173_152_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_152_6 = {3'd0, _zz_when_ArraySlice_l173_152_7};
  assign _zz_when_ArraySlice_l173_152_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_153 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_153_1);
  assign _zz_when_ArraySlice_l165_153_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_153_1 = {2'd0, _zz_when_ArraySlice_l165_153_2};
  assign _zz_when_ArraySlice_l166_153 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_153_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_153_2);
  assign _zz_when_ArraySlice_l166_153_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_153_3);
  assign _zz_when_ArraySlice_l166_153_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_153_3 = {2'd0, _zz_when_ArraySlice_l166_153_4};
  assign _zz__zz_when_ArraySlice_l112_153 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_153 = (_zz_when_ArraySlice_l113_153_1 - _zz_when_ArraySlice_l113_153_4);
  assign _zz_when_ArraySlice_l113_153_1 = (_zz_when_ArraySlice_l113_153_2 + _zz_when_ArraySlice_l113_153_3);
  assign _zz_when_ArraySlice_l113_153_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_153_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_153_4 = {1'd0, _zz_when_ArraySlice_l112_153};
  assign _zz__zz_when_ArraySlice_l173_153 = (_zz__zz_when_ArraySlice_l173_153_1 + _zz__zz_when_ArraySlice_l173_153_2);
  assign _zz__zz_when_ArraySlice_l173_153_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_153_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_153_3 = {1'd0, _zz_when_ArraySlice_l112_153};
  assign _zz_when_ArraySlice_l118_153_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_153 = _zz_when_ArraySlice_l118_153_1[5:0];
  assign _zz_when_ArraySlice_l173_153_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_153_1 = {1'd0, _zz_when_ArraySlice_l173_153_2};
  assign _zz_when_ArraySlice_l173_153_3 = (_zz_when_ArraySlice_l173_153_4 + _zz_when_ArraySlice_l173_153_9);
  assign _zz_when_ArraySlice_l173_153_4 = (_zz_when_ArraySlice_l173_153 - _zz_when_ArraySlice_l173_153_5);
  assign _zz_when_ArraySlice_l173_153_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_153_7);
  assign _zz_when_ArraySlice_l173_153_5 = {1'd0, _zz_when_ArraySlice_l173_153_6};
  assign _zz_when_ArraySlice_l173_153_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_153_7 = {2'd0, _zz_when_ArraySlice_l173_153_8};
  assign _zz_when_ArraySlice_l173_153_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_154 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_154_1);
  assign _zz_when_ArraySlice_l165_154_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_154_1 = {1'd0, _zz_when_ArraySlice_l165_154_2};
  assign _zz_when_ArraySlice_l166_154 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_154_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_154_2);
  assign _zz_when_ArraySlice_l166_154_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_154_3);
  assign _zz_when_ArraySlice_l166_154_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_154_3 = {1'd0, _zz_when_ArraySlice_l166_154_4};
  assign _zz__zz_when_ArraySlice_l112_154 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_154 = (_zz_when_ArraySlice_l113_154_1 - _zz_when_ArraySlice_l113_154_4);
  assign _zz_when_ArraySlice_l113_154_1 = (_zz_when_ArraySlice_l113_154_2 + _zz_when_ArraySlice_l113_154_3);
  assign _zz_when_ArraySlice_l113_154_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_154_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_154_4 = {1'd0, _zz_when_ArraySlice_l112_154};
  assign _zz__zz_when_ArraySlice_l173_154 = (_zz__zz_when_ArraySlice_l173_154_1 + _zz__zz_when_ArraySlice_l173_154_2);
  assign _zz__zz_when_ArraySlice_l173_154_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_154_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_154_3 = {1'd0, _zz_when_ArraySlice_l112_154};
  assign _zz_when_ArraySlice_l118_154_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_154 = _zz_when_ArraySlice_l118_154_1[5:0];
  assign _zz_when_ArraySlice_l173_154_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_154_1 = {1'd0, _zz_when_ArraySlice_l173_154_2};
  assign _zz_when_ArraySlice_l173_154_3 = (_zz_when_ArraySlice_l173_154_4 + _zz_when_ArraySlice_l173_154_9);
  assign _zz_when_ArraySlice_l173_154_4 = (_zz_when_ArraySlice_l173_154 - _zz_when_ArraySlice_l173_154_5);
  assign _zz_when_ArraySlice_l173_154_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_154_7);
  assign _zz_when_ArraySlice_l173_154_5 = {1'd0, _zz_when_ArraySlice_l173_154_6};
  assign _zz_when_ArraySlice_l173_154_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_154_7 = {1'd0, _zz_when_ArraySlice_l173_154_8};
  assign _zz_when_ArraySlice_l173_154_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_155 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_155_1);
  assign _zz_when_ArraySlice_l165_155_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_155_1 = {1'd0, _zz_when_ArraySlice_l165_155_2};
  assign _zz_when_ArraySlice_l166_155 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_155_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_155_2);
  assign _zz_when_ArraySlice_l166_155_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_155_3);
  assign _zz_when_ArraySlice_l166_155_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_155_3 = {1'd0, _zz_when_ArraySlice_l166_155_4};
  assign _zz__zz_when_ArraySlice_l112_155 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_155 = (_zz_when_ArraySlice_l113_155_1 - _zz_when_ArraySlice_l113_155_4);
  assign _zz_when_ArraySlice_l113_155_1 = (_zz_when_ArraySlice_l113_155_2 + _zz_when_ArraySlice_l113_155_3);
  assign _zz_when_ArraySlice_l113_155_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_155_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_155_4 = {1'd0, _zz_when_ArraySlice_l112_155};
  assign _zz__zz_when_ArraySlice_l173_155 = (_zz__zz_when_ArraySlice_l173_155_1 + _zz__zz_when_ArraySlice_l173_155_2);
  assign _zz__zz_when_ArraySlice_l173_155_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_155_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_155_3 = {1'd0, _zz_when_ArraySlice_l112_155};
  assign _zz_when_ArraySlice_l118_155_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_155 = _zz_when_ArraySlice_l118_155_1[5:0];
  assign _zz_when_ArraySlice_l173_155_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_155_1 = {1'd0, _zz_when_ArraySlice_l173_155_2};
  assign _zz_when_ArraySlice_l173_155_3 = (_zz_when_ArraySlice_l173_155_4 + _zz_when_ArraySlice_l173_155_9);
  assign _zz_when_ArraySlice_l173_155_4 = (_zz_when_ArraySlice_l173_155 - _zz_when_ArraySlice_l173_155_5);
  assign _zz_when_ArraySlice_l173_155_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_155_7);
  assign _zz_when_ArraySlice_l173_155_5 = {1'd0, _zz_when_ArraySlice_l173_155_6};
  assign _zz_when_ArraySlice_l173_155_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_155_7 = {1'd0, _zz_when_ArraySlice_l173_155_8};
  assign _zz_when_ArraySlice_l173_155_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_156 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_156_1);
  assign _zz_when_ArraySlice_l165_156_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_156 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_156_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_156_2);
  assign _zz_when_ArraySlice_l166_156_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_156_3);
  assign _zz_when_ArraySlice_l166_156_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_156 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_156 = (_zz_when_ArraySlice_l113_156_1 - _zz_when_ArraySlice_l113_156_4);
  assign _zz_when_ArraySlice_l113_156_1 = (_zz_when_ArraySlice_l113_156_2 + _zz_when_ArraySlice_l113_156_3);
  assign _zz_when_ArraySlice_l113_156_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_156_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_156_4 = {1'd0, _zz_when_ArraySlice_l112_156};
  assign _zz__zz_when_ArraySlice_l173_156 = (_zz__zz_when_ArraySlice_l173_156_1 + _zz__zz_when_ArraySlice_l173_156_2);
  assign _zz__zz_when_ArraySlice_l173_156_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_156_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_156_3 = {1'd0, _zz_when_ArraySlice_l112_156};
  assign _zz_when_ArraySlice_l118_156_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_156 = _zz_when_ArraySlice_l118_156_1[5:0];
  assign _zz_when_ArraySlice_l173_156_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_156_1 = {1'd0, _zz_when_ArraySlice_l173_156_2};
  assign _zz_when_ArraySlice_l173_156_3 = (_zz_when_ArraySlice_l173_156_4 + _zz_when_ArraySlice_l173_156_8);
  assign _zz_when_ArraySlice_l173_156_4 = (_zz_when_ArraySlice_l173_156 - _zz_when_ArraySlice_l173_156_5);
  assign _zz_when_ArraySlice_l173_156_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_156_7);
  assign _zz_when_ArraySlice_l173_156_5 = {1'd0, _zz_when_ArraySlice_l173_156_6};
  assign _zz_when_ArraySlice_l173_156_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_156_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_157 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_157_1);
  assign _zz_when_ArraySlice_l165_157_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_157_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_157 = {1'd0, _zz_when_ArraySlice_l166_157_1};
  assign _zz_when_ArraySlice_l166_157_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_157_3);
  assign _zz_when_ArraySlice_l166_157_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_157_4);
  assign _zz_when_ArraySlice_l166_157_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_157 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_157 = (_zz_when_ArraySlice_l113_157_1 - _zz_when_ArraySlice_l113_157_4);
  assign _zz_when_ArraySlice_l113_157_1 = (_zz_when_ArraySlice_l113_157_2 + _zz_when_ArraySlice_l113_157_3);
  assign _zz_when_ArraySlice_l113_157_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_157_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_157_4 = {1'd0, _zz_when_ArraySlice_l112_157};
  assign _zz__zz_when_ArraySlice_l173_157 = (_zz__zz_when_ArraySlice_l173_157_1 + _zz__zz_when_ArraySlice_l173_157_2);
  assign _zz__zz_when_ArraySlice_l173_157_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_157_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_157_3 = {1'd0, _zz_when_ArraySlice_l112_157};
  assign _zz_when_ArraySlice_l118_157_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_157 = _zz_when_ArraySlice_l118_157_1[5:0];
  assign _zz_when_ArraySlice_l173_157_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_157_1 = {2'd0, _zz_when_ArraySlice_l173_157_2};
  assign _zz_when_ArraySlice_l173_157_3 = (_zz_when_ArraySlice_l173_157_4 + _zz_when_ArraySlice_l173_157_8);
  assign _zz_when_ArraySlice_l173_157_4 = (_zz_when_ArraySlice_l173_157 - _zz_when_ArraySlice_l173_157_5);
  assign _zz_when_ArraySlice_l173_157_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_157_7);
  assign _zz_when_ArraySlice_l173_157_5 = {1'd0, _zz_when_ArraySlice_l173_157_6};
  assign _zz_when_ArraySlice_l173_157_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_157_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_158 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_158_1);
  assign _zz_when_ArraySlice_l165_158_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_158_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_158 = {1'd0, _zz_when_ArraySlice_l166_158_1};
  assign _zz_when_ArraySlice_l166_158_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_158_3);
  assign _zz_when_ArraySlice_l166_158_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_158_4);
  assign _zz_when_ArraySlice_l166_158_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_158 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_158 = (_zz_when_ArraySlice_l113_158_1 - _zz_when_ArraySlice_l113_158_4);
  assign _zz_when_ArraySlice_l113_158_1 = (_zz_when_ArraySlice_l113_158_2 + _zz_when_ArraySlice_l113_158_3);
  assign _zz_when_ArraySlice_l113_158_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_158_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_158_4 = {1'd0, _zz_when_ArraySlice_l112_158};
  assign _zz__zz_when_ArraySlice_l173_158 = (_zz__zz_when_ArraySlice_l173_158_1 + _zz__zz_when_ArraySlice_l173_158_2);
  assign _zz__zz_when_ArraySlice_l173_158_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_158_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_158_3 = {1'd0, _zz_when_ArraySlice_l112_158};
  assign _zz_when_ArraySlice_l118_158_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_158 = _zz_when_ArraySlice_l118_158_1[5:0];
  assign _zz_when_ArraySlice_l173_158_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_158_1 = {2'd0, _zz_when_ArraySlice_l173_158_2};
  assign _zz_when_ArraySlice_l173_158_3 = (_zz_when_ArraySlice_l173_158_4 + _zz_when_ArraySlice_l173_158_8);
  assign _zz_when_ArraySlice_l173_158_4 = (_zz_when_ArraySlice_l173_158 - _zz_when_ArraySlice_l173_158_5);
  assign _zz_when_ArraySlice_l173_158_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_158_7);
  assign _zz_when_ArraySlice_l173_158_5 = {1'd0, _zz_when_ArraySlice_l173_158_6};
  assign _zz_when_ArraySlice_l173_158_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_158_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_159 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_159_1);
  assign _zz_when_ArraySlice_l165_159_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_159_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_159 = {2'd0, _zz_when_ArraySlice_l166_159_1};
  assign _zz_when_ArraySlice_l166_159_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_159_3);
  assign _zz_when_ArraySlice_l166_159_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_159_4);
  assign _zz_when_ArraySlice_l166_159_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_159 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_159 = (_zz_when_ArraySlice_l113_159_1 - _zz_when_ArraySlice_l113_159_4);
  assign _zz_when_ArraySlice_l113_159_1 = (_zz_when_ArraySlice_l113_159_2 + _zz_when_ArraySlice_l113_159_3);
  assign _zz_when_ArraySlice_l113_159_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_159_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_159_4 = {1'd0, _zz_when_ArraySlice_l112_159};
  assign _zz__zz_when_ArraySlice_l173_159 = (_zz__zz_when_ArraySlice_l173_159_1 + _zz__zz_when_ArraySlice_l173_159_2);
  assign _zz__zz_when_ArraySlice_l173_159_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_159_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_159_3 = {1'd0, _zz_when_ArraySlice_l112_159};
  assign _zz_when_ArraySlice_l118_159_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_159 = _zz_when_ArraySlice_l118_159_1[5:0];
  assign _zz_when_ArraySlice_l173_159_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_159_1 = {3'd0, _zz_when_ArraySlice_l173_159_2};
  assign _zz_when_ArraySlice_l173_159_3 = (_zz_when_ArraySlice_l173_159_4 + _zz_when_ArraySlice_l173_159_8);
  assign _zz_when_ArraySlice_l173_159_4 = (_zz_when_ArraySlice_l173_159 - _zz_when_ArraySlice_l173_159_5);
  assign _zz_when_ArraySlice_l173_159_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_159_7);
  assign _zz_when_ArraySlice_l173_159_5 = {1'd0, _zz_when_ArraySlice_l173_159_6};
  assign _zz_when_ArraySlice_l173_159_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_159_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l401_6_1 = (_zz_when_ArraySlice_l401_6_2 + _zz_when_ArraySlice_l401_6_7);
  assign _zz_when_ArraySlice_l401_6_2 = (_zz_when_ArraySlice_l401_6_3 + _zz_when_ArraySlice_l401_6_5);
  assign _zz_when_ArraySlice_l401_6_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l401_6_4);
  assign _zz_when_ArraySlice_l401_6_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l401_6_6 = 1'b1;
  assign _zz_when_ArraySlice_l401_6_5 = {5'd0, _zz_when_ArraySlice_l401_6_6};
  assign _zz_when_ArraySlice_l401_6_7 = (bReg * 3'b110);
  assign _zz_selectReadFifo_6_15 = 1'b1;
  assign _zz_selectReadFifo_6_14 = {5'd0, _zz_selectReadFifo_6_15};
  assign _zz_when_ArraySlice_l405_6 = (_zz_when_ArraySlice_l405_6_1 % aReg);
  assign _zz_when_ArraySlice_l405_6_1 = (handshakeTimes_6_value + _zz_when_ArraySlice_l405_6_2);
  assign _zz_when_ArraySlice_l405_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l405_6_2 = {12'd0, _zz_when_ArraySlice_l405_6_3};
  assign _zz_when_ArraySlice_l409_6_1 = (selectReadFifo_6 + _zz_when_ArraySlice_l409_6_2);
  assign _zz_when_ArraySlice_l409_6_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l410_6_1 = (_zz_when_ArraySlice_l410_6_2 - _zz_when_ArraySlice_l410_6_3);
  assign _zz_when_ArraySlice_l410_6 = {7'd0, _zz_when_ArraySlice_l410_6_1};
  assign _zz_when_ArraySlice_l410_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l410_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l410_6_3 = {5'd0, _zz_when_ArraySlice_l410_6_4};
  assign _zz__zz_when_ArraySlice_l94_19 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_19 = (_zz_when_ArraySlice_l95_19_1 - _zz_when_ArraySlice_l95_19_4);
  assign _zz_when_ArraySlice_l95_19_1 = (_zz_when_ArraySlice_l95_19_2 + _zz_when_ArraySlice_l95_19_3);
  assign _zz_when_ArraySlice_l95_19_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_19_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_19_4 = {1'd0, _zz_when_ArraySlice_l94_19};
  assign _zz__zz_when_ArraySlice_l412_6 = (_zz__zz_when_ArraySlice_l412_6_1 + _zz__zz_when_ArraySlice_l412_6_2);
  assign _zz__zz_when_ArraySlice_l412_6_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l412_6_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l412_6_3 = {1'd0, _zz_when_ArraySlice_l94_19};
  assign _zz_when_ArraySlice_l99_19_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_19 = _zz_when_ArraySlice_l99_19_1[5:0];
  assign _zz_when_ArraySlice_l412_6_1 = (outSliceNumb_6_value + _zz_when_ArraySlice_l412_6_2);
  assign _zz_when_ArraySlice_l412_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l412_6_2 = {6'd0, _zz_when_ArraySlice_l412_6_3};
  assign _zz_when_ArraySlice_l412_6_4 = (_zz_when_ArraySlice_l412_6 / aReg);
  assign _zz_selectReadFifo_6_16 = (selectReadFifo_6 - _zz_selectReadFifo_6_17);
  assign _zz_selectReadFifo_6_17 = {3'd0, bReg};
  assign _zz_selectReadFifo_6_19 = 1'b1;
  assign _zz_selectReadFifo_6_18 = {5'd0, _zz_selectReadFifo_6_19};
  assign _zz_selectReadFifo_6_20 = (selectReadFifo_6 + _zz_selectReadFifo_6_21);
  assign _zz_selectReadFifo_6_21 = (3'b111 * bReg);
  assign _zz_selectReadFifo_6_23 = 1'b1;
  assign _zz_selectReadFifo_6_22 = {5'd0, _zz_selectReadFifo_6_23};
  assign _zz_when_ArraySlice_l165_160 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_160_1);
  assign _zz_when_ArraySlice_l165_160_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_160_1 = {3'd0, _zz_when_ArraySlice_l165_160_2};
  assign _zz_when_ArraySlice_l166_160 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_160_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_160_3);
  assign _zz_when_ArraySlice_l166_160_1 = {1'd0, _zz_when_ArraySlice_l166_160_2};
  assign _zz_when_ArraySlice_l166_160_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_160_4);
  assign _zz_when_ArraySlice_l166_160_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_160_4 = {3'd0, _zz_when_ArraySlice_l166_160_5};
  assign _zz__zz_when_ArraySlice_l112_160 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_160 = (_zz_when_ArraySlice_l113_160_1 - _zz_when_ArraySlice_l113_160_4);
  assign _zz_when_ArraySlice_l113_160_1 = (_zz_when_ArraySlice_l113_160_2 + _zz_when_ArraySlice_l113_160_3);
  assign _zz_when_ArraySlice_l113_160_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_160_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_160_4 = {1'd0, _zz_when_ArraySlice_l112_160};
  assign _zz__zz_when_ArraySlice_l173_160 = (_zz__zz_when_ArraySlice_l173_160_1 + _zz__zz_when_ArraySlice_l173_160_2);
  assign _zz__zz_when_ArraySlice_l173_160_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_160_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_160_3 = {1'd0, _zz_when_ArraySlice_l112_160};
  assign _zz_when_ArraySlice_l118_160_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_160 = _zz_when_ArraySlice_l118_160_1[5:0];
  assign _zz_when_ArraySlice_l173_160_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_160_2 = (_zz_when_ArraySlice_l173_160_3 + _zz_when_ArraySlice_l173_160_8);
  assign _zz_when_ArraySlice_l173_160_3 = (_zz_when_ArraySlice_l173_160 - _zz_when_ArraySlice_l173_160_4);
  assign _zz_when_ArraySlice_l173_160_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_160_6);
  assign _zz_when_ArraySlice_l173_160_4 = {1'd0, _zz_when_ArraySlice_l173_160_5};
  assign _zz_when_ArraySlice_l173_160_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_160_6 = {3'd0, _zz_when_ArraySlice_l173_160_7};
  assign _zz_when_ArraySlice_l173_160_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_161 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_161_1);
  assign _zz_when_ArraySlice_l165_161_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_161_1 = {2'd0, _zz_when_ArraySlice_l165_161_2};
  assign _zz_when_ArraySlice_l166_161 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_161_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_161_2);
  assign _zz_when_ArraySlice_l166_161_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_161_3);
  assign _zz_when_ArraySlice_l166_161_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_161_3 = {2'd0, _zz_when_ArraySlice_l166_161_4};
  assign _zz__zz_when_ArraySlice_l112_161 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_161 = (_zz_when_ArraySlice_l113_161_1 - _zz_when_ArraySlice_l113_161_4);
  assign _zz_when_ArraySlice_l113_161_1 = (_zz_when_ArraySlice_l113_161_2 + _zz_when_ArraySlice_l113_161_3);
  assign _zz_when_ArraySlice_l113_161_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_161_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_161_4 = {1'd0, _zz_when_ArraySlice_l112_161};
  assign _zz__zz_when_ArraySlice_l173_161 = (_zz__zz_when_ArraySlice_l173_161_1 + _zz__zz_when_ArraySlice_l173_161_2);
  assign _zz__zz_when_ArraySlice_l173_161_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_161_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_161_3 = {1'd0, _zz_when_ArraySlice_l112_161};
  assign _zz_when_ArraySlice_l118_161_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_161 = _zz_when_ArraySlice_l118_161_1[5:0];
  assign _zz_when_ArraySlice_l173_161_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_161_1 = {1'd0, _zz_when_ArraySlice_l173_161_2};
  assign _zz_when_ArraySlice_l173_161_3 = (_zz_when_ArraySlice_l173_161_4 + _zz_when_ArraySlice_l173_161_9);
  assign _zz_when_ArraySlice_l173_161_4 = (_zz_when_ArraySlice_l173_161 - _zz_when_ArraySlice_l173_161_5);
  assign _zz_when_ArraySlice_l173_161_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_161_7);
  assign _zz_when_ArraySlice_l173_161_5 = {1'd0, _zz_when_ArraySlice_l173_161_6};
  assign _zz_when_ArraySlice_l173_161_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_161_7 = {2'd0, _zz_when_ArraySlice_l173_161_8};
  assign _zz_when_ArraySlice_l173_161_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_162 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_162_1);
  assign _zz_when_ArraySlice_l165_162_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_162_1 = {1'd0, _zz_when_ArraySlice_l165_162_2};
  assign _zz_when_ArraySlice_l166_162 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_162_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_162_2);
  assign _zz_when_ArraySlice_l166_162_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_162_3);
  assign _zz_when_ArraySlice_l166_162_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_162_3 = {1'd0, _zz_when_ArraySlice_l166_162_4};
  assign _zz__zz_when_ArraySlice_l112_162 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_162 = (_zz_when_ArraySlice_l113_162_1 - _zz_when_ArraySlice_l113_162_4);
  assign _zz_when_ArraySlice_l113_162_1 = (_zz_when_ArraySlice_l113_162_2 + _zz_when_ArraySlice_l113_162_3);
  assign _zz_when_ArraySlice_l113_162_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_162_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_162_4 = {1'd0, _zz_when_ArraySlice_l112_162};
  assign _zz__zz_when_ArraySlice_l173_162 = (_zz__zz_when_ArraySlice_l173_162_1 + _zz__zz_when_ArraySlice_l173_162_2);
  assign _zz__zz_when_ArraySlice_l173_162_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_162_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_162_3 = {1'd0, _zz_when_ArraySlice_l112_162};
  assign _zz_when_ArraySlice_l118_162_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_162 = _zz_when_ArraySlice_l118_162_1[5:0];
  assign _zz_when_ArraySlice_l173_162_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_162_1 = {1'd0, _zz_when_ArraySlice_l173_162_2};
  assign _zz_when_ArraySlice_l173_162_3 = (_zz_when_ArraySlice_l173_162_4 + _zz_when_ArraySlice_l173_162_9);
  assign _zz_when_ArraySlice_l173_162_4 = (_zz_when_ArraySlice_l173_162 - _zz_when_ArraySlice_l173_162_5);
  assign _zz_when_ArraySlice_l173_162_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_162_7);
  assign _zz_when_ArraySlice_l173_162_5 = {1'd0, _zz_when_ArraySlice_l173_162_6};
  assign _zz_when_ArraySlice_l173_162_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_162_7 = {1'd0, _zz_when_ArraySlice_l173_162_8};
  assign _zz_when_ArraySlice_l173_162_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_163 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_163_1);
  assign _zz_when_ArraySlice_l165_163_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_163_1 = {1'd0, _zz_when_ArraySlice_l165_163_2};
  assign _zz_when_ArraySlice_l166_163 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_163_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_163_2);
  assign _zz_when_ArraySlice_l166_163_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_163_3);
  assign _zz_when_ArraySlice_l166_163_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_163_3 = {1'd0, _zz_when_ArraySlice_l166_163_4};
  assign _zz__zz_when_ArraySlice_l112_163 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_163 = (_zz_when_ArraySlice_l113_163_1 - _zz_when_ArraySlice_l113_163_4);
  assign _zz_when_ArraySlice_l113_163_1 = (_zz_when_ArraySlice_l113_163_2 + _zz_when_ArraySlice_l113_163_3);
  assign _zz_when_ArraySlice_l113_163_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_163_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_163_4 = {1'd0, _zz_when_ArraySlice_l112_163};
  assign _zz__zz_when_ArraySlice_l173_163 = (_zz__zz_when_ArraySlice_l173_163_1 + _zz__zz_when_ArraySlice_l173_163_2);
  assign _zz__zz_when_ArraySlice_l173_163_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_163_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_163_3 = {1'd0, _zz_when_ArraySlice_l112_163};
  assign _zz_when_ArraySlice_l118_163_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_163 = _zz_when_ArraySlice_l118_163_1[5:0];
  assign _zz_when_ArraySlice_l173_163_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_163_1 = {1'd0, _zz_when_ArraySlice_l173_163_2};
  assign _zz_when_ArraySlice_l173_163_3 = (_zz_when_ArraySlice_l173_163_4 + _zz_when_ArraySlice_l173_163_9);
  assign _zz_when_ArraySlice_l173_163_4 = (_zz_when_ArraySlice_l173_163 - _zz_when_ArraySlice_l173_163_5);
  assign _zz_when_ArraySlice_l173_163_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_163_7);
  assign _zz_when_ArraySlice_l173_163_5 = {1'd0, _zz_when_ArraySlice_l173_163_6};
  assign _zz_when_ArraySlice_l173_163_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_163_7 = {1'd0, _zz_when_ArraySlice_l173_163_8};
  assign _zz_when_ArraySlice_l173_163_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_164 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_164_1);
  assign _zz_when_ArraySlice_l165_164_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_164 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_164_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_164_2);
  assign _zz_when_ArraySlice_l166_164_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_164_3);
  assign _zz_when_ArraySlice_l166_164_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_164 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_164 = (_zz_when_ArraySlice_l113_164_1 - _zz_when_ArraySlice_l113_164_4);
  assign _zz_when_ArraySlice_l113_164_1 = (_zz_when_ArraySlice_l113_164_2 + _zz_when_ArraySlice_l113_164_3);
  assign _zz_when_ArraySlice_l113_164_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_164_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_164_4 = {1'd0, _zz_when_ArraySlice_l112_164};
  assign _zz__zz_when_ArraySlice_l173_164 = (_zz__zz_when_ArraySlice_l173_164_1 + _zz__zz_when_ArraySlice_l173_164_2);
  assign _zz__zz_when_ArraySlice_l173_164_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_164_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_164_3 = {1'd0, _zz_when_ArraySlice_l112_164};
  assign _zz_when_ArraySlice_l118_164_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_164 = _zz_when_ArraySlice_l118_164_1[5:0];
  assign _zz_when_ArraySlice_l173_164_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_164_1 = {1'd0, _zz_when_ArraySlice_l173_164_2};
  assign _zz_when_ArraySlice_l173_164_3 = (_zz_when_ArraySlice_l173_164_4 + _zz_when_ArraySlice_l173_164_8);
  assign _zz_when_ArraySlice_l173_164_4 = (_zz_when_ArraySlice_l173_164 - _zz_when_ArraySlice_l173_164_5);
  assign _zz_when_ArraySlice_l173_164_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_164_7);
  assign _zz_when_ArraySlice_l173_164_5 = {1'd0, _zz_when_ArraySlice_l173_164_6};
  assign _zz_when_ArraySlice_l173_164_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_164_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_165 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_165_1);
  assign _zz_when_ArraySlice_l165_165_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_165_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_165 = {1'd0, _zz_when_ArraySlice_l166_165_1};
  assign _zz_when_ArraySlice_l166_165_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_165_3);
  assign _zz_when_ArraySlice_l166_165_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_165_4);
  assign _zz_when_ArraySlice_l166_165_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_165 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_165 = (_zz_when_ArraySlice_l113_165_1 - _zz_when_ArraySlice_l113_165_4);
  assign _zz_when_ArraySlice_l113_165_1 = (_zz_when_ArraySlice_l113_165_2 + _zz_when_ArraySlice_l113_165_3);
  assign _zz_when_ArraySlice_l113_165_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_165_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_165_4 = {1'd0, _zz_when_ArraySlice_l112_165};
  assign _zz__zz_when_ArraySlice_l173_165 = (_zz__zz_when_ArraySlice_l173_165_1 + _zz__zz_when_ArraySlice_l173_165_2);
  assign _zz__zz_when_ArraySlice_l173_165_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_165_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_165_3 = {1'd0, _zz_when_ArraySlice_l112_165};
  assign _zz_when_ArraySlice_l118_165_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_165 = _zz_when_ArraySlice_l118_165_1[5:0];
  assign _zz_when_ArraySlice_l173_165_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_165_1 = {2'd0, _zz_when_ArraySlice_l173_165_2};
  assign _zz_when_ArraySlice_l173_165_3 = (_zz_when_ArraySlice_l173_165_4 + _zz_when_ArraySlice_l173_165_8);
  assign _zz_when_ArraySlice_l173_165_4 = (_zz_when_ArraySlice_l173_165 - _zz_when_ArraySlice_l173_165_5);
  assign _zz_when_ArraySlice_l173_165_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_165_7);
  assign _zz_when_ArraySlice_l173_165_5 = {1'd0, _zz_when_ArraySlice_l173_165_6};
  assign _zz_when_ArraySlice_l173_165_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_165_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_166 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_166_1);
  assign _zz_when_ArraySlice_l165_166_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_166_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_166 = {1'd0, _zz_when_ArraySlice_l166_166_1};
  assign _zz_when_ArraySlice_l166_166_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_166_3);
  assign _zz_when_ArraySlice_l166_166_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_166_4);
  assign _zz_when_ArraySlice_l166_166_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_166 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_166 = (_zz_when_ArraySlice_l113_166_1 - _zz_when_ArraySlice_l113_166_4);
  assign _zz_when_ArraySlice_l113_166_1 = (_zz_when_ArraySlice_l113_166_2 + _zz_when_ArraySlice_l113_166_3);
  assign _zz_when_ArraySlice_l113_166_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_166_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_166_4 = {1'd0, _zz_when_ArraySlice_l112_166};
  assign _zz__zz_when_ArraySlice_l173_166 = (_zz__zz_when_ArraySlice_l173_166_1 + _zz__zz_when_ArraySlice_l173_166_2);
  assign _zz__zz_when_ArraySlice_l173_166_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_166_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_166_3 = {1'd0, _zz_when_ArraySlice_l112_166};
  assign _zz_when_ArraySlice_l118_166_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_166 = _zz_when_ArraySlice_l118_166_1[5:0];
  assign _zz_when_ArraySlice_l173_166_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_166_1 = {2'd0, _zz_when_ArraySlice_l173_166_2};
  assign _zz_when_ArraySlice_l173_166_3 = (_zz_when_ArraySlice_l173_166_4 + _zz_when_ArraySlice_l173_166_8);
  assign _zz_when_ArraySlice_l173_166_4 = (_zz_when_ArraySlice_l173_166 - _zz_when_ArraySlice_l173_166_5);
  assign _zz_when_ArraySlice_l173_166_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_166_7);
  assign _zz_when_ArraySlice_l173_166_5 = {1'd0, _zz_when_ArraySlice_l173_166_6};
  assign _zz_when_ArraySlice_l173_166_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_166_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_167 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_167_1);
  assign _zz_when_ArraySlice_l165_167_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_167_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_167 = {2'd0, _zz_when_ArraySlice_l166_167_1};
  assign _zz_when_ArraySlice_l166_167_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_167_3);
  assign _zz_when_ArraySlice_l166_167_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_167_4);
  assign _zz_when_ArraySlice_l166_167_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_167 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_167 = (_zz_when_ArraySlice_l113_167_1 - _zz_when_ArraySlice_l113_167_4);
  assign _zz_when_ArraySlice_l113_167_1 = (_zz_when_ArraySlice_l113_167_2 + _zz_when_ArraySlice_l113_167_3);
  assign _zz_when_ArraySlice_l113_167_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_167_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_167_4 = {1'd0, _zz_when_ArraySlice_l112_167};
  assign _zz__zz_when_ArraySlice_l173_167 = (_zz__zz_when_ArraySlice_l173_167_1 + _zz__zz_when_ArraySlice_l173_167_2);
  assign _zz__zz_when_ArraySlice_l173_167_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_167_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_167_3 = {1'd0, _zz_when_ArraySlice_l112_167};
  assign _zz_when_ArraySlice_l118_167_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_167 = _zz_when_ArraySlice_l118_167_1[5:0];
  assign _zz_when_ArraySlice_l173_167_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_167_1 = {3'd0, _zz_when_ArraySlice_l173_167_2};
  assign _zz_when_ArraySlice_l173_167_3 = (_zz_when_ArraySlice_l173_167_4 + _zz_when_ArraySlice_l173_167_8);
  assign _zz_when_ArraySlice_l173_167_4 = (_zz_when_ArraySlice_l173_167 - _zz_when_ArraySlice_l173_167_5);
  assign _zz_when_ArraySlice_l173_167_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_167_7);
  assign _zz_when_ArraySlice_l173_167_5 = {1'd0, _zz_when_ArraySlice_l173_167_6};
  assign _zz_when_ArraySlice_l173_167_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_167_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l421_6_1 = (_zz_when_ArraySlice_l421_6_2 + _zz_when_ArraySlice_l421_6_7);
  assign _zz_when_ArraySlice_l421_6_2 = (_zz_when_ArraySlice_l421_6_3 + _zz_when_ArraySlice_l421_6_5);
  assign _zz_when_ArraySlice_l421_6_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l421_6_4);
  assign _zz_when_ArraySlice_l421_6_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l421_6_6 = 1'b1;
  assign _zz_when_ArraySlice_l421_6_5 = {5'd0, _zz_when_ArraySlice_l421_6_6};
  assign _zz_when_ArraySlice_l421_6_7 = (bReg * 3'b110);
  assign _zz_selectReadFifo_6_25 = 1'b1;
  assign _zz_selectReadFifo_6_24 = {5'd0, _zz_selectReadFifo_6_25};
  assign _zz_when_ArraySlice_l425_6 = (_zz_when_ArraySlice_l425_6_1 % aReg);
  assign _zz_when_ArraySlice_l425_6_1 = (handshakeTimes_6_value + _zz_when_ArraySlice_l425_6_2);
  assign _zz_when_ArraySlice_l425_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l425_6_2 = {12'd0, _zz_when_ArraySlice_l425_6_3};
  assign _zz_when_ArraySlice_l436_6_1 = (_zz_when_ArraySlice_l436_6_2 - _zz_when_ArraySlice_l436_6_3);
  assign _zz_when_ArraySlice_l436_6 = {7'd0, _zz_when_ArraySlice_l436_6_1};
  assign _zz_when_ArraySlice_l436_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l436_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l436_6_3 = {5'd0, _zz_when_ArraySlice_l436_6_4};
  assign _zz__zz_when_ArraySlice_l94_20 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_20 = (_zz_when_ArraySlice_l95_20_1 - _zz_when_ArraySlice_l95_20_4);
  assign _zz_when_ArraySlice_l95_20_1 = (_zz_when_ArraySlice_l95_20_2 + _zz_when_ArraySlice_l95_20_3);
  assign _zz_when_ArraySlice_l95_20_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_20_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_20_4 = {1'd0, _zz_when_ArraySlice_l94_20};
  assign _zz__zz_when_ArraySlice_l437_6 = (_zz__zz_when_ArraySlice_l437_6_1 + _zz__zz_when_ArraySlice_l437_6_2);
  assign _zz__zz_when_ArraySlice_l437_6_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l437_6_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l437_6_3 = {1'd0, _zz_when_ArraySlice_l94_20};
  assign _zz_when_ArraySlice_l99_20_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_20 = _zz_when_ArraySlice_l99_20_1[5:0];
  assign _zz_when_ArraySlice_l437_6_1 = (outSliceNumb_6_value + _zz_when_ArraySlice_l437_6_2);
  assign _zz_when_ArraySlice_l437_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l437_6_2 = {6'd0, _zz_when_ArraySlice_l437_6_3};
  assign _zz_when_ArraySlice_l437_6_4 = (_zz_when_ArraySlice_l437_6 / aReg);
  assign _zz_selectReadFifo_6_26 = (selectReadFifo_6 - _zz_selectReadFifo_6_27);
  assign _zz_selectReadFifo_6_27 = {3'd0, bReg};
  assign _zz_selectReadFifo_6_29 = 1'b1;
  assign _zz_selectReadFifo_6_28 = {5'd0, _zz_selectReadFifo_6_29};
  assign _zz_when_ArraySlice_l165_168 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_168_1);
  assign _zz_when_ArraySlice_l165_168_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_168_1 = {3'd0, _zz_when_ArraySlice_l165_168_2};
  assign _zz_when_ArraySlice_l166_168 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_168_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_168_3);
  assign _zz_when_ArraySlice_l166_168_1 = {1'd0, _zz_when_ArraySlice_l166_168_2};
  assign _zz_when_ArraySlice_l166_168_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_168_4);
  assign _zz_when_ArraySlice_l166_168_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_168_4 = {3'd0, _zz_when_ArraySlice_l166_168_5};
  assign _zz__zz_when_ArraySlice_l112_168 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_168 = (_zz_when_ArraySlice_l113_168_1 - _zz_when_ArraySlice_l113_168_4);
  assign _zz_when_ArraySlice_l113_168_1 = (_zz_when_ArraySlice_l113_168_2 + _zz_when_ArraySlice_l113_168_3);
  assign _zz_when_ArraySlice_l113_168_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_168_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_168_4 = {1'd0, _zz_when_ArraySlice_l112_168};
  assign _zz__zz_when_ArraySlice_l173_168 = (_zz__zz_when_ArraySlice_l173_168_1 + _zz__zz_when_ArraySlice_l173_168_2);
  assign _zz__zz_when_ArraySlice_l173_168_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_168_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_168_3 = {1'd0, _zz_when_ArraySlice_l112_168};
  assign _zz_when_ArraySlice_l118_168_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_168 = _zz_when_ArraySlice_l118_168_1[5:0];
  assign _zz_when_ArraySlice_l173_168_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_168_2 = (_zz_when_ArraySlice_l173_168_3 + _zz_when_ArraySlice_l173_168_8);
  assign _zz_when_ArraySlice_l173_168_3 = (_zz_when_ArraySlice_l173_168 - _zz_when_ArraySlice_l173_168_4);
  assign _zz_when_ArraySlice_l173_168_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_168_6);
  assign _zz_when_ArraySlice_l173_168_4 = {1'd0, _zz_when_ArraySlice_l173_168_5};
  assign _zz_when_ArraySlice_l173_168_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_168_6 = {3'd0, _zz_when_ArraySlice_l173_168_7};
  assign _zz_when_ArraySlice_l173_168_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_169 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_169_1);
  assign _zz_when_ArraySlice_l165_169_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_169_1 = {2'd0, _zz_when_ArraySlice_l165_169_2};
  assign _zz_when_ArraySlice_l166_169 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_169_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_169_2);
  assign _zz_when_ArraySlice_l166_169_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_169_3);
  assign _zz_when_ArraySlice_l166_169_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_169_3 = {2'd0, _zz_when_ArraySlice_l166_169_4};
  assign _zz__zz_when_ArraySlice_l112_169 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_169 = (_zz_when_ArraySlice_l113_169_1 - _zz_when_ArraySlice_l113_169_4);
  assign _zz_when_ArraySlice_l113_169_1 = (_zz_when_ArraySlice_l113_169_2 + _zz_when_ArraySlice_l113_169_3);
  assign _zz_when_ArraySlice_l113_169_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_169_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_169_4 = {1'd0, _zz_when_ArraySlice_l112_169};
  assign _zz__zz_when_ArraySlice_l173_169 = (_zz__zz_when_ArraySlice_l173_169_1 + _zz__zz_when_ArraySlice_l173_169_2);
  assign _zz__zz_when_ArraySlice_l173_169_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_169_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_169_3 = {1'd0, _zz_when_ArraySlice_l112_169};
  assign _zz_when_ArraySlice_l118_169_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_169 = _zz_when_ArraySlice_l118_169_1[5:0];
  assign _zz_when_ArraySlice_l173_169_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_169_1 = {1'd0, _zz_when_ArraySlice_l173_169_2};
  assign _zz_when_ArraySlice_l173_169_3 = (_zz_when_ArraySlice_l173_169_4 + _zz_when_ArraySlice_l173_169_9);
  assign _zz_when_ArraySlice_l173_169_4 = (_zz_when_ArraySlice_l173_169 - _zz_when_ArraySlice_l173_169_5);
  assign _zz_when_ArraySlice_l173_169_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_169_7);
  assign _zz_when_ArraySlice_l173_169_5 = {1'd0, _zz_when_ArraySlice_l173_169_6};
  assign _zz_when_ArraySlice_l173_169_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_169_7 = {2'd0, _zz_when_ArraySlice_l173_169_8};
  assign _zz_when_ArraySlice_l173_169_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_170 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_170_1);
  assign _zz_when_ArraySlice_l165_170_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_170_1 = {1'd0, _zz_when_ArraySlice_l165_170_2};
  assign _zz_when_ArraySlice_l166_170 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_170_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_170_2);
  assign _zz_when_ArraySlice_l166_170_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_170_3);
  assign _zz_when_ArraySlice_l166_170_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_170_3 = {1'd0, _zz_when_ArraySlice_l166_170_4};
  assign _zz__zz_when_ArraySlice_l112_170 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_170 = (_zz_when_ArraySlice_l113_170_1 - _zz_when_ArraySlice_l113_170_4);
  assign _zz_when_ArraySlice_l113_170_1 = (_zz_when_ArraySlice_l113_170_2 + _zz_when_ArraySlice_l113_170_3);
  assign _zz_when_ArraySlice_l113_170_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_170_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_170_4 = {1'd0, _zz_when_ArraySlice_l112_170};
  assign _zz__zz_when_ArraySlice_l173_170 = (_zz__zz_when_ArraySlice_l173_170_1 + _zz__zz_when_ArraySlice_l173_170_2);
  assign _zz__zz_when_ArraySlice_l173_170_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_170_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_170_3 = {1'd0, _zz_when_ArraySlice_l112_170};
  assign _zz_when_ArraySlice_l118_170_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_170 = _zz_when_ArraySlice_l118_170_1[5:0];
  assign _zz_when_ArraySlice_l173_170_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_170_1 = {1'd0, _zz_when_ArraySlice_l173_170_2};
  assign _zz_when_ArraySlice_l173_170_3 = (_zz_when_ArraySlice_l173_170_4 + _zz_when_ArraySlice_l173_170_9);
  assign _zz_when_ArraySlice_l173_170_4 = (_zz_when_ArraySlice_l173_170 - _zz_when_ArraySlice_l173_170_5);
  assign _zz_when_ArraySlice_l173_170_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_170_7);
  assign _zz_when_ArraySlice_l173_170_5 = {1'd0, _zz_when_ArraySlice_l173_170_6};
  assign _zz_when_ArraySlice_l173_170_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_170_7 = {1'd0, _zz_when_ArraySlice_l173_170_8};
  assign _zz_when_ArraySlice_l173_170_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_171 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_171_1);
  assign _zz_when_ArraySlice_l165_171_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_171_1 = {1'd0, _zz_when_ArraySlice_l165_171_2};
  assign _zz_when_ArraySlice_l166_171 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_171_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_171_2);
  assign _zz_when_ArraySlice_l166_171_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_171_3);
  assign _zz_when_ArraySlice_l166_171_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_171_3 = {1'd0, _zz_when_ArraySlice_l166_171_4};
  assign _zz__zz_when_ArraySlice_l112_171 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_171 = (_zz_when_ArraySlice_l113_171_1 - _zz_when_ArraySlice_l113_171_4);
  assign _zz_when_ArraySlice_l113_171_1 = (_zz_when_ArraySlice_l113_171_2 + _zz_when_ArraySlice_l113_171_3);
  assign _zz_when_ArraySlice_l113_171_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_171_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_171_4 = {1'd0, _zz_when_ArraySlice_l112_171};
  assign _zz__zz_when_ArraySlice_l173_171 = (_zz__zz_when_ArraySlice_l173_171_1 + _zz__zz_when_ArraySlice_l173_171_2);
  assign _zz__zz_when_ArraySlice_l173_171_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_171_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_171_3 = {1'd0, _zz_when_ArraySlice_l112_171};
  assign _zz_when_ArraySlice_l118_171_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_171 = _zz_when_ArraySlice_l118_171_1[5:0];
  assign _zz_when_ArraySlice_l173_171_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_171_1 = {1'd0, _zz_when_ArraySlice_l173_171_2};
  assign _zz_when_ArraySlice_l173_171_3 = (_zz_when_ArraySlice_l173_171_4 + _zz_when_ArraySlice_l173_171_9);
  assign _zz_when_ArraySlice_l173_171_4 = (_zz_when_ArraySlice_l173_171 - _zz_when_ArraySlice_l173_171_5);
  assign _zz_when_ArraySlice_l173_171_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_171_7);
  assign _zz_when_ArraySlice_l173_171_5 = {1'd0, _zz_when_ArraySlice_l173_171_6};
  assign _zz_when_ArraySlice_l173_171_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_171_7 = {1'd0, _zz_when_ArraySlice_l173_171_8};
  assign _zz_when_ArraySlice_l173_171_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_172 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_172_1);
  assign _zz_when_ArraySlice_l165_172_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_172 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_172_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_172_2);
  assign _zz_when_ArraySlice_l166_172_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_172_3);
  assign _zz_when_ArraySlice_l166_172_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_172 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_172 = (_zz_when_ArraySlice_l113_172_1 - _zz_when_ArraySlice_l113_172_4);
  assign _zz_when_ArraySlice_l113_172_1 = (_zz_when_ArraySlice_l113_172_2 + _zz_when_ArraySlice_l113_172_3);
  assign _zz_when_ArraySlice_l113_172_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_172_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_172_4 = {1'd0, _zz_when_ArraySlice_l112_172};
  assign _zz__zz_when_ArraySlice_l173_172 = (_zz__zz_when_ArraySlice_l173_172_1 + _zz__zz_when_ArraySlice_l173_172_2);
  assign _zz__zz_when_ArraySlice_l173_172_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_172_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_172_3 = {1'd0, _zz_when_ArraySlice_l112_172};
  assign _zz_when_ArraySlice_l118_172_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_172 = _zz_when_ArraySlice_l118_172_1[5:0];
  assign _zz_when_ArraySlice_l173_172_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_172_1 = {1'd0, _zz_when_ArraySlice_l173_172_2};
  assign _zz_when_ArraySlice_l173_172_3 = (_zz_when_ArraySlice_l173_172_4 + _zz_when_ArraySlice_l173_172_8);
  assign _zz_when_ArraySlice_l173_172_4 = (_zz_when_ArraySlice_l173_172 - _zz_when_ArraySlice_l173_172_5);
  assign _zz_when_ArraySlice_l173_172_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_172_7);
  assign _zz_when_ArraySlice_l173_172_5 = {1'd0, _zz_when_ArraySlice_l173_172_6};
  assign _zz_when_ArraySlice_l173_172_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_172_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_173 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_173_1);
  assign _zz_when_ArraySlice_l165_173_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_173_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_173 = {1'd0, _zz_when_ArraySlice_l166_173_1};
  assign _zz_when_ArraySlice_l166_173_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_173_3);
  assign _zz_when_ArraySlice_l166_173_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_173_4);
  assign _zz_when_ArraySlice_l166_173_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_173 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_173 = (_zz_when_ArraySlice_l113_173_1 - _zz_when_ArraySlice_l113_173_4);
  assign _zz_when_ArraySlice_l113_173_1 = (_zz_when_ArraySlice_l113_173_2 + _zz_when_ArraySlice_l113_173_3);
  assign _zz_when_ArraySlice_l113_173_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_173_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_173_4 = {1'd0, _zz_when_ArraySlice_l112_173};
  assign _zz__zz_when_ArraySlice_l173_173 = (_zz__zz_when_ArraySlice_l173_173_1 + _zz__zz_when_ArraySlice_l173_173_2);
  assign _zz__zz_when_ArraySlice_l173_173_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_173_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_173_3 = {1'd0, _zz_when_ArraySlice_l112_173};
  assign _zz_when_ArraySlice_l118_173_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_173 = _zz_when_ArraySlice_l118_173_1[5:0];
  assign _zz_when_ArraySlice_l173_173_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_173_1 = {2'd0, _zz_when_ArraySlice_l173_173_2};
  assign _zz_when_ArraySlice_l173_173_3 = (_zz_when_ArraySlice_l173_173_4 + _zz_when_ArraySlice_l173_173_8);
  assign _zz_when_ArraySlice_l173_173_4 = (_zz_when_ArraySlice_l173_173 - _zz_when_ArraySlice_l173_173_5);
  assign _zz_when_ArraySlice_l173_173_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_173_7);
  assign _zz_when_ArraySlice_l173_173_5 = {1'd0, _zz_when_ArraySlice_l173_173_6};
  assign _zz_when_ArraySlice_l173_173_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_173_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_174 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_174_1);
  assign _zz_when_ArraySlice_l165_174_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_174_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_174 = {1'd0, _zz_when_ArraySlice_l166_174_1};
  assign _zz_when_ArraySlice_l166_174_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_174_3);
  assign _zz_when_ArraySlice_l166_174_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_174_4);
  assign _zz_when_ArraySlice_l166_174_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_174 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_174 = (_zz_when_ArraySlice_l113_174_1 - _zz_when_ArraySlice_l113_174_4);
  assign _zz_when_ArraySlice_l113_174_1 = (_zz_when_ArraySlice_l113_174_2 + _zz_when_ArraySlice_l113_174_3);
  assign _zz_when_ArraySlice_l113_174_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_174_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_174_4 = {1'd0, _zz_when_ArraySlice_l112_174};
  assign _zz__zz_when_ArraySlice_l173_174 = (_zz__zz_when_ArraySlice_l173_174_1 + _zz__zz_when_ArraySlice_l173_174_2);
  assign _zz__zz_when_ArraySlice_l173_174_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_174_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_174_3 = {1'd0, _zz_when_ArraySlice_l112_174};
  assign _zz_when_ArraySlice_l118_174_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_174 = _zz_when_ArraySlice_l118_174_1[5:0];
  assign _zz_when_ArraySlice_l173_174_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_174_1 = {2'd0, _zz_when_ArraySlice_l173_174_2};
  assign _zz_when_ArraySlice_l173_174_3 = (_zz_when_ArraySlice_l173_174_4 + _zz_when_ArraySlice_l173_174_8);
  assign _zz_when_ArraySlice_l173_174_4 = (_zz_when_ArraySlice_l173_174 - _zz_when_ArraySlice_l173_174_5);
  assign _zz_when_ArraySlice_l173_174_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_174_7);
  assign _zz_when_ArraySlice_l173_174_5 = {1'd0, _zz_when_ArraySlice_l173_174_6};
  assign _zz_when_ArraySlice_l173_174_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_174_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_175 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_175_1);
  assign _zz_when_ArraySlice_l165_175_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_175_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_175 = {2'd0, _zz_when_ArraySlice_l166_175_1};
  assign _zz_when_ArraySlice_l166_175_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_175_3);
  assign _zz_when_ArraySlice_l166_175_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_175_4);
  assign _zz_when_ArraySlice_l166_175_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_175 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_175 = (_zz_when_ArraySlice_l113_175_1 - _zz_when_ArraySlice_l113_175_4);
  assign _zz_when_ArraySlice_l113_175_1 = (_zz_when_ArraySlice_l113_175_2 + _zz_when_ArraySlice_l113_175_3);
  assign _zz_when_ArraySlice_l113_175_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_175_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_175_4 = {1'd0, _zz_when_ArraySlice_l112_175};
  assign _zz__zz_when_ArraySlice_l173_175 = (_zz__zz_when_ArraySlice_l173_175_1 + _zz__zz_when_ArraySlice_l173_175_2);
  assign _zz__zz_when_ArraySlice_l173_175_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_175_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_175_3 = {1'd0, _zz_when_ArraySlice_l112_175};
  assign _zz_when_ArraySlice_l118_175_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_175 = _zz_when_ArraySlice_l118_175_1[5:0];
  assign _zz_when_ArraySlice_l173_175_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_175_1 = {3'd0, _zz_when_ArraySlice_l173_175_2};
  assign _zz_when_ArraySlice_l173_175_3 = (_zz_when_ArraySlice_l173_175_4 + _zz_when_ArraySlice_l173_175_8);
  assign _zz_when_ArraySlice_l173_175_4 = (_zz_when_ArraySlice_l173_175 - _zz_when_ArraySlice_l173_175_5);
  assign _zz_when_ArraySlice_l173_175_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_175_7);
  assign _zz_when_ArraySlice_l173_175_5 = {1'd0, _zz_when_ArraySlice_l173_175_6};
  assign _zz_when_ArraySlice_l173_175_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_175_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_6_31 = 1'b1;
  assign _zz_selectReadFifo_6_30 = {5'd0, _zz_selectReadFifo_6_31};
  assign _zz_when_ArraySlice_l448_6 = (_zz_when_ArraySlice_l448_6_1 % aReg);
  assign _zz_when_ArraySlice_l448_6_1 = (handshakeTimes_6_value + _zz_when_ArraySlice_l448_6_2);
  assign _zz_when_ArraySlice_l448_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l448_6_2 = {12'd0, _zz_when_ArraySlice_l448_6_3};
  assign _zz_when_ArraySlice_l434_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l434_6_1);
  assign _zz_when_ArraySlice_l434_6_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l455_6_1 = (_zz_when_ArraySlice_l455_6_2 - _zz_when_ArraySlice_l455_6_3);
  assign _zz_when_ArraySlice_l455_6 = {7'd0, _zz_when_ArraySlice_l455_6_1};
  assign _zz_when_ArraySlice_l455_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l455_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l455_6_3 = {5'd0, _zz_when_ArraySlice_l455_6_4};
  assign _zz_when_ArraySlice_l373_7 = (selectReadFifo_7 + _zz_when_ArraySlice_l373_7_1);
  assign _zz_when_ArraySlice_l373_7_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l374_7_1 = (selectReadFifo_7 + _zz_when_ArraySlice_l374_7_2);
  assign _zz_when_ArraySlice_l374_7_2 = (bReg * 3'b111);
  assign _zz__zz_outputStreamArrayData_7_valid = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l380_7_1 = 1'b1;
  assign _zz_when_ArraySlice_l380_7 = {6'd0, _zz_when_ArraySlice_l380_7_1};
  assign _zz_when_ArraySlice_l380_7_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l380_7_4);
  assign _zz_when_ArraySlice_l380_7_4 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l381_7_1 = (_zz_when_ArraySlice_l381_7_2 - _zz_when_ArraySlice_l381_7_3);
  assign _zz_when_ArraySlice_l381_7 = {7'd0, _zz_when_ArraySlice_l381_7_1};
  assign _zz_when_ArraySlice_l381_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l381_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l381_7_3 = {5'd0, _zz_when_ArraySlice_l381_7_4};
  assign _zz_selectReadFifo_7 = (selectReadFifo_7 - _zz_selectReadFifo_7_1);
  assign _zz_selectReadFifo_7_1 = {3'd0, bReg};
  assign _zz_selectReadFifo_7_3 = 1'b1;
  assign _zz_selectReadFifo_7_2 = {5'd0, _zz_selectReadFifo_7_3};
  assign _zz_selectReadFifo_7_5 = 1'b1;
  assign _zz_selectReadFifo_7_4 = {5'd0, _zz_selectReadFifo_7_5};
  assign _zz_when_ArraySlice_l384_7 = (_zz_when_ArraySlice_l384_7_1 % aReg);
  assign _zz_when_ArraySlice_l384_7_1 = (handshakeTimes_7_value + _zz_when_ArraySlice_l384_7_2);
  assign _zz_when_ArraySlice_l384_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l384_7_2 = {12'd0, _zz_when_ArraySlice_l384_7_3};
  assign _zz_when_ArraySlice_l389_7_1 = (selectReadFifo_7 + _zz_when_ArraySlice_l389_7_2);
  assign _zz_when_ArraySlice_l389_7_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l389_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l389_7_3 = {6'd0, _zz_when_ArraySlice_l389_7_4};
  assign _zz_when_ArraySlice_l390_7_1 = (_zz_when_ArraySlice_l390_7_2 - _zz_when_ArraySlice_l390_7_3);
  assign _zz_when_ArraySlice_l390_7 = {7'd0, _zz_when_ArraySlice_l390_7_1};
  assign _zz_when_ArraySlice_l390_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l390_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l390_7_3 = {5'd0, _zz_when_ArraySlice_l390_7_4};
  assign _zz__zz_when_ArraySlice_l94_21 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_21 = (_zz_when_ArraySlice_l95_21_1 - _zz_when_ArraySlice_l95_21_4);
  assign _zz_when_ArraySlice_l95_21_1 = (_zz_when_ArraySlice_l95_21_2 + _zz_when_ArraySlice_l95_21_3);
  assign _zz_when_ArraySlice_l95_21_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_21_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_21_4 = {1'd0, _zz_when_ArraySlice_l94_21};
  assign _zz__zz_when_ArraySlice_l392_7 = (_zz__zz_when_ArraySlice_l392_7_1 + _zz__zz_when_ArraySlice_l392_7_2);
  assign _zz__zz_when_ArraySlice_l392_7_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l392_7_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l392_7_3 = {1'd0, _zz_when_ArraySlice_l94_21};
  assign _zz_when_ArraySlice_l99_21_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_21 = _zz_when_ArraySlice_l99_21_1[5:0];
  assign _zz_when_ArraySlice_l392_7_1 = (outSliceNumb_7_value + _zz_when_ArraySlice_l392_7_2);
  assign _zz_when_ArraySlice_l392_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l392_7_2 = {6'd0, _zz_when_ArraySlice_l392_7_3};
  assign _zz_when_ArraySlice_l392_7_4 = (_zz_when_ArraySlice_l392_7 / aReg);
  assign _zz_selectReadFifo_7_6 = (selectReadFifo_7 - _zz_selectReadFifo_7_7);
  assign _zz_selectReadFifo_7_7 = {3'd0, bReg};
  assign _zz_selectReadFifo_7_9 = 1'b1;
  assign _zz_selectReadFifo_7_8 = {5'd0, _zz_selectReadFifo_7_9};
  assign _zz_selectReadFifo_7_10 = (selectReadFifo_7 + _zz_selectReadFifo_7_11);
  assign _zz_selectReadFifo_7_11 = (3'b111 * bReg);
  assign _zz_selectReadFifo_7_13 = 1'b1;
  assign _zz_selectReadFifo_7_12 = {5'd0, _zz_selectReadFifo_7_13};
  assign _zz_when_ArraySlice_l165_176 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_176_1);
  assign _zz_when_ArraySlice_l165_176_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_176_1 = {3'd0, _zz_when_ArraySlice_l165_176_2};
  assign _zz_when_ArraySlice_l166_176 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_176_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_176_3);
  assign _zz_when_ArraySlice_l166_176_1 = {1'd0, _zz_when_ArraySlice_l166_176_2};
  assign _zz_when_ArraySlice_l166_176_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_176_4);
  assign _zz_when_ArraySlice_l166_176_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_176_4 = {3'd0, _zz_when_ArraySlice_l166_176_5};
  assign _zz__zz_when_ArraySlice_l112_176 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_176 = (_zz_when_ArraySlice_l113_176_1 - _zz_when_ArraySlice_l113_176_4);
  assign _zz_when_ArraySlice_l113_176_1 = (_zz_when_ArraySlice_l113_176_2 + _zz_when_ArraySlice_l113_176_3);
  assign _zz_when_ArraySlice_l113_176_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_176_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_176_4 = {1'd0, _zz_when_ArraySlice_l112_176};
  assign _zz__zz_when_ArraySlice_l173_176 = (_zz__zz_when_ArraySlice_l173_176_1 + _zz__zz_when_ArraySlice_l173_176_2);
  assign _zz__zz_when_ArraySlice_l173_176_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_176_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_176_3 = {1'd0, _zz_when_ArraySlice_l112_176};
  assign _zz_when_ArraySlice_l118_176_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_176 = _zz_when_ArraySlice_l118_176_1[5:0];
  assign _zz_when_ArraySlice_l173_176_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_176_2 = (_zz_when_ArraySlice_l173_176_3 + _zz_when_ArraySlice_l173_176_8);
  assign _zz_when_ArraySlice_l173_176_3 = (_zz_when_ArraySlice_l173_176 - _zz_when_ArraySlice_l173_176_4);
  assign _zz_when_ArraySlice_l173_176_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_176_6);
  assign _zz_when_ArraySlice_l173_176_4 = {1'd0, _zz_when_ArraySlice_l173_176_5};
  assign _zz_when_ArraySlice_l173_176_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_176_6 = {3'd0, _zz_when_ArraySlice_l173_176_7};
  assign _zz_when_ArraySlice_l173_176_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_177 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_177_1);
  assign _zz_when_ArraySlice_l165_177_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_177_1 = {2'd0, _zz_when_ArraySlice_l165_177_2};
  assign _zz_when_ArraySlice_l166_177 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_177_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_177_2);
  assign _zz_when_ArraySlice_l166_177_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_177_3);
  assign _zz_when_ArraySlice_l166_177_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_177_3 = {2'd0, _zz_when_ArraySlice_l166_177_4};
  assign _zz__zz_when_ArraySlice_l112_177 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_177 = (_zz_when_ArraySlice_l113_177_1 - _zz_when_ArraySlice_l113_177_4);
  assign _zz_when_ArraySlice_l113_177_1 = (_zz_when_ArraySlice_l113_177_2 + _zz_when_ArraySlice_l113_177_3);
  assign _zz_when_ArraySlice_l113_177_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_177_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_177_4 = {1'd0, _zz_when_ArraySlice_l112_177};
  assign _zz__zz_when_ArraySlice_l173_177 = (_zz__zz_when_ArraySlice_l173_177_1 + _zz__zz_when_ArraySlice_l173_177_2);
  assign _zz__zz_when_ArraySlice_l173_177_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_177_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_177_3 = {1'd0, _zz_when_ArraySlice_l112_177};
  assign _zz_when_ArraySlice_l118_177_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_177 = _zz_when_ArraySlice_l118_177_1[5:0];
  assign _zz_when_ArraySlice_l173_177_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_177_1 = {1'd0, _zz_when_ArraySlice_l173_177_2};
  assign _zz_when_ArraySlice_l173_177_3 = (_zz_when_ArraySlice_l173_177_4 + _zz_when_ArraySlice_l173_177_9);
  assign _zz_when_ArraySlice_l173_177_4 = (_zz_when_ArraySlice_l173_177 - _zz_when_ArraySlice_l173_177_5);
  assign _zz_when_ArraySlice_l173_177_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_177_7);
  assign _zz_when_ArraySlice_l173_177_5 = {1'd0, _zz_when_ArraySlice_l173_177_6};
  assign _zz_when_ArraySlice_l173_177_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_177_7 = {2'd0, _zz_when_ArraySlice_l173_177_8};
  assign _zz_when_ArraySlice_l173_177_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_178 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_178_1);
  assign _zz_when_ArraySlice_l165_178_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_178_1 = {1'd0, _zz_when_ArraySlice_l165_178_2};
  assign _zz_when_ArraySlice_l166_178 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_178_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_178_2);
  assign _zz_when_ArraySlice_l166_178_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_178_3);
  assign _zz_when_ArraySlice_l166_178_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_178_3 = {1'd0, _zz_when_ArraySlice_l166_178_4};
  assign _zz__zz_when_ArraySlice_l112_178 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_178 = (_zz_when_ArraySlice_l113_178_1 - _zz_when_ArraySlice_l113_178_4);
  assign _zz_when_ArraySlice_l113_178_1 = (_zz_when_ArraySlice_l113_178_2 + _zz_when_ArraySlice_l113_178_3);
  assign _zz_when_ArraySlice_l113_178_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_178_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_178_4 = {1'd0, _zz_when_ArraySlice_l112_178};
  assign _zz__zz_when_ArraySlice_l173_178 = (_zz__zz_when_ArraySlice_l173_178_1 + _zz__zz_when_ArraySlice_l173_178_2);
  assign _zz__zz_when_ArraySlice_l173_178_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_178_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_178_3 = {1'd0, _zz_when_ArraySlice_l112_178};
  assign _zz_when_ArraySlice_l118_178_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_178 = _zz_when_ArraySlice_l118_178_1[5:0];
  assign _zz_when_ArraySlice_l173_178_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_178_1 = {1'd0, _zz_when_ArraySlice_l173_178_2};
  assign _zz_when_ArraySlice_l173_178_3 = (_zz_when_ArraySlice_l173_178_4 + _zz_when_ArraySlice_l173_178_9);
  assign _zz_when_ArraySlice_l173_178_4 = (_zz_when_ArraySlice_l173_178 - _zz_when_ArraySlice_l173_178_5);
  assign _zz_when_ArraySlice_l173_178_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_178_7);
  assign _zz_when_ArraySlice_l173_178_5 = {1'd0, _zz_when_ArraySlice_l173_178_6};
  assign _zz_when_ArraySlice_l173_178_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_178_7 = {1'd0, _zz_when_ArraySlice_l173_178_8};
  assign _zz_when_ArraySlice_l173_178_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_179 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_179_1);
  assign _zz_when_ArraySlice_l165_179_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_179_1 = {1'd0, _zz_when_ArraySlice_l165_179_2};
  assign _zz_when_ArraySlice_l166_179 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_179_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_179_2);
  assign _zz_when_ArraySlice_l166_179_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_179_3);
  assign _zz_when_ArraySlice_l166_179_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_179_3 = {1'd0, _zz_when_ArraySlice_l166_179_4};
  assign _zz__zz_when_ArraySlice_l112_179 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_179 = (_zz_when_ArraySlice_l113_179_1 - _zz_when_ArraySlice_l113_179_4);
  assign _zz_when_ArraySlice_l113_179_1 = (_zz_when_ArraySlice_l113_179_2 + _zz_when_ArraySlice_l113_179_3);
  assign _zz_when_ArraySlice_l113_179_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_179_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_179_4 = {1'd0, _zz_when_ArraySlice_l112_179};
  assign _zz__zz_when_ArraySlice_l173_179 = (_zz__zz_when_ArraySlice_l173_179_1 + _zz__zz_when_ArraySlice_l173_179_2);
  assign _zz__zz_when_ArraySlice_l173_179_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_179_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_179_3 = {1'd0, _zz_when_ArraySlice_l112_179};
  assign _zz_when_ArraySlice_l118_179_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_179 = _zz_when_ArraySlice_l118_179_1[5:0];
  assign _zz_when_ArraySlice_l173_179_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_179_1 = {1'd0, _zz_when_ArraySlice_l173_179_2};
  assign _zz_when_ArraySlice_l173_179_3 = (_zz_when_ArraySlice_l173_179_4 + _zz_when_ArraySlice_l173_179_9);
  assign _zz_when_ArraySlice_l173_179_4 = (_zz_when_ArraySlice_l173_179 - _zz_when_ArraySlice_l173_179_5);
  assign _zz_when_ArraySlice_l173_179_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_179_7);
  assign _zz_when_ArraySlice_l173_179_5 = {1'd0, _zz_when_ArraySlice_l173_179_6};
  assign _zz_when_ArraySlice_l173_179_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_179_7 = {1'd0, _zz_when_ArraySlice_l173_179_8};
  assign _zz_when_ArraySlice_l173_179_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_180 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_180_1);
  assign _zz_when_ArraySlice_l165_180_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_180 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_180_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_180_2);
  assign _zz_when_ArraySlice_l166_180_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_180_3);
  assign _zz_when_ArraySlice_l166_180_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_180 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_180 = (_zz_when_ArraySlice_l113_180_1 - _zz_when_ArraySlice_l113_180_4);
  assign _zz_when_ArraySlice_l113_180_1 = (_zz_when_ArraySlice_l113_180_2 + _zz_when_ArraySlice_l113_180_3);
  assign _zz_when_ArraySlice_l113_180_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_180_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_180_4 = {1'd0, _zz_when_ArraySlice_l112_180};
  assign _zz__zz_when_ArraySlice_l173_180 = (_zz__zz_when_ArraySlice_l173_180_1 + _zz__zz_when_ArraySlice_l173_180_2);
  assign _zz__zz_when_ArraySlice_l173_180_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_180_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_180_3 = {1'd0, _zz_when_ArraySlice_l112_180};
  assign _zz_when_ArraySlice_l118_180_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_180 = _zz_when_ArraySlice_l118_180_1[5:0];
  assign _zz_when_ArraySlice_l173_180_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_180_1 = {1'd0, _zz_when_ArraySlice_l173_180_2};
  assign _zz_when_ArraySlice_l173_180_3 = (_zz_when_ArraySlice_l173_180_4 + _zz_when_ArraySlice_l173_180_8);
  assign _zz_when_ArraySlice_l173_180_4 = (_zz_when_ArraySlice_l173_180 - _zz_when_ArraySlice_l173_180_5);
  assign _zz_when_ArraySlice_l173_180_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_180_7);
  assign _zz_when_ArraySlice_l173_180_5 = {1'd0, _zz_when_ArraySlice_l173_180_6};
  assign _zz_when_ArraySlice_l173_180_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_180_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_181 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_181_1);
  assign _zz_when_ArraySlice_l165_181_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_181_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_181 = {1'd0, _zz_when_ArraySlice_l166_181_1};
  assign _zz_when_ArraySlice_l166_181_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_181_3);
  assign _zz_when_ArraySlice_l166_181_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_181_4);
  assign _zz_when_ArraySlice_l166_181_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_181 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_181 = (_zz_when_ArraySlice_l113_181_1 - _zz_when_ArraySlice_l113_181_4);
  assign _zz_when_ArraySlice_l113_181_1 = (_zz_when_ArraySlice_l113_181_2 + _zz_when_ArraySlice_l113_181_3);
  assign _zz_when_ArraySlice_l113_181_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_181_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_181_4 = {1'd0, _zz_when_ArraySlice_l112_181};
  assign _zz__zz_when_ArraySlice_l173_181 = (_zz__zz_when_ArraySlice_l173_181_1 + _zz__zz_when_ArraySlice_l173_181_2);
  assign _zz__zz_when_ArraySlice_l173_181_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_181_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_181_3 = {1'd0, _zz_when_ArraySlice_l112_181};
  assign _zz_when_ArraySlice_l118_181_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_181 = _zz_when_ArraySlice_l118_181_1[5:0];
  assign _zz_when_ArraySlice_l173_181_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_181_1 = {2'd0, _zz_when_ArraySlice_l173_181_2};
  assign _zz_when_ArraySlice_l173_181_3 = (_zz_when_ArraySlice_l173_181_4 + _zz_when_ArraySlice_l173_181_8);
  assign _zz_when_ArraySlice_l173_181_4 = (_zz_when_ArraySlice_l173_181 - _zz_when_ArraySlice_l173_181_5);
  assign _zz_when_ArraySlice_l173_181_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_181_7);
  assign _zz_when_ArraySlice_l173_181_5 = {1'd0, _zz_when_ArraySlice_l173_181_6};
  assign _zz_when_ArraySlice_l173_181_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_181_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_182 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_182_1);
  assign _zz_when_ArraySlice_l165_182_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_182_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_182 = {1'd0, _zz_when_ArraySlice_l166_182_1};
  assign _zz_when_ArraySlice_l166_182_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_182_3);
  assign _zz_when_ArraySlice_l166_182_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_182_4);
  assign _zz_when_ArraySlice_l166_182_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_182 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_182 = (_zz_when_ArraySlice_l113_182_1 - _zz_when_ArraySlice_l113_182_4);
  assign _zz_when_ArraySlice_l113_182_1 = (_zz_when_ArraySlice_l113_182_2 + _zz_when_ArraySlice_l113_182_3);
  assign _zz_when_ArraySlice_l113_182_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_182_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_182_4 = {1'd0, _zz_when_ArraySlice_l112_182};
  assign _zz__zz_when_ArraySlice_l173_182 = (_zz__zz_when_ArraySlice_l173_182_1 + _zz__zz_when_ArraySlice_l173_182_2);
  assign _zz__zz_when_ArraySlice_l173_182_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_182_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_182_3 = {1'd0, _zz_when_ArraySlice_l112_182};
  assign _zz_when_ArraySlice_l118_182_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_182 = _zz_when_ArraySlice_l118_182_1[5:0];
  assign _zz_when_ArraySlice_l173_182_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_182_1 = {2'd0, _zz_when_ArraySlice_l173_182_2};
  assign _zz_when_ArraySlice_l173_182_3 = (_zz_when_ArraySlice_l173_182_4 + _zz_when_ArraySlice_l173_182_8);
  assign _zz_when_ArraySlice_l173_182_4 = (_zz_when_ArraySlice_l173_182 - _zz_when_ArraySlice_l173_182_5);
  assign _zz_when_ArraySlice_l173_182_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_182_7);
  assign _zz_when_ArraySlice_l173_182_5 = {1'd0, _zz_when_ArraySlice_l173_182_6};
  assign _zz_when_ArraySlice_l173_182_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_182_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_183 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_183_1);
  assign _zz_when_ArraySlice_l165_183_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_183_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_183 = {2'd0, _zz_when_ArraySlice_l166_183_1};
  assign _zz_when_ArraySlice_l166_183_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_183_3);
  assign _zz_when_ArraySlice_l166_183_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_183_4);
  assign _zz_when_ArraySlice_l166_183_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_183 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_183 = (_zz_when_ArraySlice_l113_183_1 - _zz_when_ArraySlice_l113_183_4);
  assign _zz_when_ArraySlice_l113_183_1 = (_zz_when_ArraySlice_l113_183_2 + _zz_when_ArraySlice_l113_183_3);
  assign _zz_when_ArraySlice_l113_183_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_183_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_183_4 = {1'd0, _zz_when_ArraySlice_l112_183};
  assign _zz__zz_when_ArraySlice_l173_183 = (_zz__zz_when_ArraySlice_l173_183_1 + _zz__zz_when_ArraySlice_l173_183_2);
  assign _zz__zz_when_ArraySlice_l173_183_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_183_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_183_3 = {1'd0, _zz_when_ArraySlice_l112_183};
  assign _zz_when_ArraySlice_l118_183_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_183 = _zz_when_ArraySlice_l118_183_1[5:0];
  assign _zz_when_ArraySlice_l173_183_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_183_1 = {3'd0, _zz_when_ArraySlice_l173_183_2};
  assign _zz_when_ArraySlice_l173_183_3 = (_zz_when_ArraySlice_l173_183_4 + _zz_when_ArraySlice_l173_183_8);
  assign _zz_when_ArraySlice_l173_183_4 = (_zz_when_ArraySlice_l173_183 - _zz_when_ArraySlice_l173_183_5);
  assign _zz_when_ArraySlice_l173_183_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_183_7);
  assign _zz_when_ArraySlice_l173_183_5 = {1'd0, _zz_when_ArraySlice_l173_183_6};
  assign _zz_when_ArraySlice_l173_183_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_183_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l401_7_1 = (_zz_when_ArraySlice_l401_7_2 + _zz_when_ArraySlice_l401_7_7);
  assign _zz_when_ArraySlice_l401_7_2 = (_zz_when_ArraySlice_l401_7_3 + _zz_when_ArraySlice_l401_7_5);
  assign _zz_when_ArraySlice_l401_7_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l401_7_4);
  assign _zz_when_ArraySlice_l401_7_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l401_7_6 = 1'b1;
  assign _zz_when_ArraySlice_l401_7_5 = {5'd0, _zz_when_ArraySlice_l401_7_6};
  assign _zz_when_ArraySlice_l401_7_7 = (bReg * 3'b111);
  assign _zz_selectReadFifo_7_15 = 1'b1;
  assign _zz_selectReadFifo_7_14 = {5'd0, _zz_selectReadFifo_7_15};
  assign _zz_when_ArraySlice_l405_7 = (_zz_when_ArraySlice_l405_7_1 % aReg);
  assign _zz_when_ArraySlice_l405_7_1 = (handshakeTimes_7_value + _zz_when_ArraySlice_l405_7_2);
  assign _zz_when_ArraySlice_l405_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l405_7_2 = {12'd0, _zz_when_ArraySlice_l405_7_3};
  assign _zz_when_ArraySlice_l409_7_1 = (selectReadFifo_7 + _zz_when_ArraySlice_l409_7_2);
  assign _zz_when_ArraySlice_l409_7_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l410_7_1 = (_zz_when_ArraySlice_l410_7_2 - _zz_when_ArraySlice_l410_7_3);
  assign _zz_when_ArraySlice_l410_7 = {7'd0, _zz_when_ArraySlice_l410_7_1};
  assign _zz_when_ArraySlice_l410_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l410_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l410_7_3 = {5'd0, _zz_when_ArraySlice_l410_7_4};
  assign _zz__zz_when_ArraySlice_l94_22 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_22 = (_zz_when_ArraySlice_l95_22_1 - _zz_when_ArraySlice_l95_22_4);
  assign _zz_when_ArraySlice_l95_22_1 = (_zz_when_ArraySlice_l95_22_2 + _zz_when_ArraySlice_l95_22_3);
  assign _zz_when_ArraySlice_l95_22_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_22_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_22_4 = {1'd0, _zz_when_ArraySlice_l94_22};
  assign _zz__zz_when_ArraySlice_l412_7 = (_zz__zz_when_ArraySlice_l412_7_1 + _zz__zz_when_ArraySlice_l412_7_2);
  assign _zz__zz_when_ArraySlice_l412_7_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l412_7_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l412_7_3 = {1'd0, _zz_when_ArraySlice_l94_22};
  assign _zz_when_ArraySlice_l99_22_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_22 = _zz_when_ArraySlice_l99_22_1[5:0];
  assign _zz_when_ArraySlice_l412_7_1 = (outSliceNumb_7_value + _zz_when_ArraySlice_l412_7_2);
  assign _zz_when_ArraySlice_l412_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l412_7_2 = {6'd0, _zz_when_ArraySlice_l412_7_3};
  assign _zz_when_ArraySlice_l412_7_4 = (_zz_when_ArraySlice_l412_7 / aReg);
  assign _zz_selectReadFifo_7_16 = (selectReadFifo_7 - _zz_selectReadFifo_7_17);
  assign _zz_selectReadFifo_7_17 = {3'd0, bReg};
  assign _zz_selectReadFifo_7_19 = 1'b1;
  assign _zz_selectReadFifo_7_18 = {5'd0, _zz_selectReadFifo_7_19};
  assign _zz_selectReadFifo_7_20 = (selectReadFifo_7 + _zz_selectReadFifo_7_21);
  assign _zz_selectReadFifo_7_21 = (3'b111 * bReg);
  assign _zz_selectReadFifo_7_23 = 1'b1;
  assign _zz_selectReadFifo_7_22 = {5'd0, _zz_selectReadFifo_7_23};
  assign _zz_when_ArraySlice_l165_184 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_184_1);
  assign _zz_when_ArraySlice_l165_184_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_184_1 = {3'd0, _zz_when_ArraySlice_l165_184_2};
  assign _zz_when_ArraySlice_l166_184 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_184_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_184_3);
  assign _zz_when_ArraySlice_l166_184_1 = {1'd0, _zz_when_ArraySlice_l166_184_2};
  assign _zz_when_ArraySlice_l166_184_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_184_4);
  assign _zz_when_ArraySlice_l166_184_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_184_4 = {3'd0, _zz_when_ArraySlice_l166_184_5};
  assign _zz__zz_when_ArraySlice_l112_184 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_184 = (_zz_when_ArraySlice_l113_184_1 - _zz_when_ArraySlice_l113_184_4);
  assign _zz_when_ArraySlice_l113_184_1 = (_zz_when_ArraySlice_l113_184_2 + _zz_when_ArraySlice_l113_184_3);
  assign _zz_when_ArraySlice_l113_184_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_184_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_184_4 = {1'd0, _zz_when_ArraySlice_l112_184};
  assign _zz__zz_when_ArraySlice_l173_184 = (_zz__zz_when_ArraySlice_l173_184_1 + _zz__zz_when_ArraySlice_l173_184_2);
  assign _zz__zz_when_ArraySlice_l173_184_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_184_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_184_3 = {1'd0, _zz_when_ArraySlice_l112_184};
  assign _zz_when_ArraySlice_l118_184_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_184 = _zz_when_ArraySlice_l118_184_1[5:0];
  assign _zz_when_ArraySlice_l173_184_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_184_2 = (_zz_when_ArraySlice_l173_184_3 + _zz_when_ArraySlice_l173_184_8);
  assign _zz_when_ArraySlice_l173_184_3 = (_zz_when_ArraySlice_l173_184 - _zz_when_ArraySlice_l173_184_4);
  assign _zz_when_ArraySlice_l173_184_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_184_6);
  assign _zz_when_ArraySlice_l173_184_4 = {1'd0, _zz_when_ArraySlice_l173_184_5};
  assign _zz_when_ArraySlice_l173_184_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_184_6 = {3'd0, _zz_when_ArraySlice_l173_184_7};
  assign _zz_when_ArraySlice_l173_184_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_185 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_185_1);
  assign _zz_when_ArraySlice_l165_185_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_185_1 = {2'd0, _zz_when_ArraySlice_l165_185_2};
  assign _zz_when_ArraySlice_l166_185 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_185_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_185_2);
  assign _zz_when_ArraySlice_l166_185_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_185_3);
  assign _zz_when_ArraySlice_l166_185_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_185_3 = {2'd0, _zz_when_ArraySlice_l166_185_4};
  assign _zz__zz_when_ArraySlice_l112_185 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_185 = (_zz_when_ArraySlice_l113_185_1 - _zz_when_ArraySlice_l113_185_4);
  assign _zz_when_ArraySlice_l113_185_1 = (_zz_when_ArraySlice_l113_185_2 + _zz_when_ArraySlice_l113_185_3);
  assign _zz_when_ArraySlice_l113_185_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_185_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_185_4 = {1'd0, _zz_when_ArraySlice_l112_185};
  assign _zz__zz_when_ArraySlice_l173_185 = (_zz__zz_when_ArraySlice_l173_185_1 + _zz__zz_when_ArraySlice_l173_185_2);
  assign _zz__zz_when_ArraySlice_l173_185_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_185_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_185_3 = {1'd0, _zz_when_ArraySlice_l112_185};
  assign _zz_when_ArraySlice_l118_185_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_185 = _zz_when_ArraySlice_l118_185_1[5:0];
  assign _zz_when_ArraySlice_l173_185_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_185_1 = {1'd0, _zz_when_ArraySlice_l173_185_2};
  assign _zz_when_ArraySlice_l173_185_3 = (_zz_when_ArraySlice_l173_185_4 + _zz_when_ArraySlice_l173_185_9);
  assign _zz_when_ArraySlice_l173_185_4 = (_zz_when_ArraySlice_l173_185 - _zz_when_ArraySlice_l173_185_5);
  assign _zz_when_ArraySlice_l173_185_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_185_7);
  assign _zz_when_ArraySlice_l173_185_5 = {1'd0, _zz_when_ArraySlice_l173_185_6};
  assign _zz_when_ArraySlice_l173_185_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_185_7 = {2'd0, _zz_when_ArraySlice_l173_185_8};
  assign _zz_when_ArraySlice_l173_185_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_186 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_186_1);
  assign _zz_when_ArraySlice_l165_186_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_186_1 = {1'd0, _zz_when_ArraySlice_l165_186_2};
  assign _zz_when_ArraySlice_l166_186 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_186_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_186_2);
  assign _zz_when_ArraySlice_l166_186_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_186_3);
  assign _zz_when_ArraySlice_l166_186_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_186_3 = {1'd0, _zz_when_ArraySlice_l166_186_4};
  assign _zz__zz_when_ArraySlice_l112_186 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_186 = (_zz_when_ArraySlice_l113_186_1 - _zz_when_ArraySlice_l113_186_4);
  assign _zz_when_ArraySlice_l113_186_1 = (_zz_when_ArraySlice_l113_186_2 + _zz_when_ArraySlice_l113_186_3);
  assign _zz_when_ArraySlice_l113_186_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_186_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_186_4 = {1'd0, _zz_when_ArraySlice_l112_186};
  assign _zz__zz_when_ArraySlice_l173_186 = (_zz__zz_when_ArraySlice_l173_186_1 + _zz__zz_when_ArraySlice_l173_186_2);
  assign _zz__zz_when_ArraySlice_l173_186_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_186_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_186_3 = {1'd0, _zz_when_ArraySlice_l112_186};
  assign _zz_when_ArraySlice_l118_186_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_186 = _zz_when_ArraySlice_l118_186_1[5:0];
  assign _zz_when_ArraySlice_l173_186_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_186_1 = {1'd0, _zz_when_ArraySlice_l173_186_2};
  assign _zz_when_ArraySlice_l173_186_3 = (_zz_when_ArraySlice_l173_186_4 + _zz_when_ArraySlice_l173_186_9);
  assign _zz_when_ArraySlice_l173_186_4 = (_zz_when_ArraySlice_l173_186 - _zz_when_ArraySlice_l173_186_5);
  assign _zz_when_ArraySlice_l173_186_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_186_7);
  assign _zz_when_ArraySlice_l173_186_5 = {1'd0, _zz_when_ArraySlice_l173_186_6};
  assign _zz_when_ArraySlice_l173_186_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_186_7 = {1'd0, _zz_when_ArraySlice_l173_186_8};
  assign _zz_when_ArraySlice_l173_186_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_187 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_187_1);
  assign _zz_when_ArraySlice_l165_187_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_187_1 = {1'd0, _zz_when_ArraySlice_l165_187_2};
  assign _zz_when_ArraySlice_l166_187 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_187_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_187_2);
  assign _zz_when_ArraySlice_l166_187_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_187_3);
  assign _zz_when_ArraySlice_l166_187_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_187_3 = {1'd0, _zz_when_ArraySlice_l166_187_4};
  assign _zz__zz_when_ArraySlice_l112_187 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_187 = (_zz_when_ArraySlice_l113_187_1 - _zz_when_ArraySlice_l113_187_4);
  assign _zz_when_ArraySlice_l113_187_1 = (_zz_when_ArraySlice_l113_187_2 + _zz_when_ArraySlice_l113_187_3);
  assign _zz_when_ArraySlice_l113_187_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_187_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_187_4 = {1'd0, _zz_when_ArraySlice_l112_187};
  assign _zz__zz_when_ArraySlice_l173_187 = (_zz__zz_when_ArraySlice_l173_187_1 + _zz__zz_when_ArraySlice_l173_187_2);
  assign _zz__zz_when_ArraySlice_l173_187_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_187_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_187_3 = {1'd0, _zz_when_ArraySlice_l112_187};
  assign _zz_when_ArraySlice_l118_187_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_187 = _zz_when_ArraySlice_l118_187_1[5:0];
  assign _zz_when_ArraySlice_l173_187_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_187_1 = {1'd0, _zz_when_ArraySlice_l173_187_2};
  assign _zz_when_ArraySlice_l173_187_3 = (_zz_when_ArraySlice_l173_187_4 + _zz_when_ArraySlice_l173_187_9);
  assign _zz_when_ArraySlice_l173_187_4 = (_zz_when_ArraySlice_l173_187 - _zz_when_ArraySlice_l173_187_5);
  assign _zz_when_ArraySlice_l173_187_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_187_7);
  assign _zz_when_ArraySlice_l173_187_5 = {1'd0, _zz_when_ArraySlice_l173_187_6};
  assign _zz_when_ArraySlice_l173_187_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_187_7 = {1'd0, _zz_when_ArraySlice_l173_187_8};
  assign _zz_when_ArraySlice_l173_187_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_188 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_188_1);
  assign _zz_when_ArraySlice_l165_188_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_188 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_188_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_188_2);
  assign _zz_when_ArraySlice_l166_188_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_188_3);
  assign _zz_when_ArraySlice_l166_188_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_188 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_188 = (_zz_when_ArraySlice_l113_188_1 - _zz_when_ArraySlice_l113_188_4);
  assign _zz_when_ArraySlice_l113_188_1 = (_zz_when_ArraySlice_l113_188_2 + _zz_when_ArraySlice_l113_188_3);
  assign _zz_when_ArraySlice_l113_188_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_188_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_188_4 = {1'd0, _zz_when_ArraySlice_l112_188};
  assign _zz__zz_when_ArraySlice_l173_188 = (_zz__zz_when_ArraySlice_l173_188_1 + _zz__zz_when_ArraySlice_l173_188_2);
  assign _zz__zz_when_ArraySlice_l173_188_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_188_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_188_3 = {1'd0, _zz_when_ArraySlice_l112_188};
  assign _zz_when_ArraySlice_l118_188_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_188 = _zz_when_ArraySlice_l118_188_1[5:0];
  assign _zz_when_ArraySlice_l173_188_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_188_1 = {1'd0, _zz_when_ArraySlice_l173_188_2};
  assign _zz_when_ArraySlice_l173_188_3 = (_zz_when_ArraySlice_l173_188_4 + _zz_when_ArraySlice_l173_188_8);
  assign _zz_when_ArraySlice_l173_188_4 = (_zz_when_ArraySlice_l173_188 - _zz_when_ArraySlice_l173_188_5);
  assign _zz_when_ArraySlice_l173_188_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_188_7);
  assign _zz_when_ArraySlice_l173_188_5 = {1'd0, _zz_when_ArraySlice_l173_188_6};
  assign _zz_when_ArraySlice_l173_188_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_188_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_189 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_189_1);
  assign _zz_when_ArraySlice_l165_189_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_189_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_189 = {1'd0, _zz_when_ArraySlice_l166_189_1};
  assign _zz_when_ArraySlice_l166_189_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_189_3);
  assign _zz_when_ArraySlice_l166_189_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_189_4);
  assign _zz_when_ArraySlice_l166_189_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_189 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_189 = (_zz_when_ArraySlice_l113_189_1 - _zz_when_ArraySlice_l113_189_4);
  assign _zz_when_ArraySlice_l113_189_1 = (_zz_when_ArraySlice_l113_189_2 + _zz_when_ArraySlice_l113_189_3);
  assign _zz_when_ArraySlice_l113_189_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_189_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_189_4 = {1'd0, _zz_when_ArraySlice_l112_189};
  assign _zz__zz_when_ArraySlice_l173_189 = (_zz__zz_when_ArraySlice_l173_189_1 + _zz__zz_when_ArraySlice_l173_189_2);
  assign _zz__zz_when_ArraySlice_l173_189_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_189_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_189_3 = {1'd0, _zz_when_ArraySlice_l112_189};
  assign _zz_when_ArraySlice_l118_189_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_189 = _zz_when_ArraySlice_l118_189_1[5:0];
  assign _zz_when_ArraySlice_l173_189_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_189_1 = {2'd0, _zz_when_ArraySlice_l173_189_2};
  assign _zz_when_ArraySlice_l173_189_3 = (_zz_when_ArraySlice_l173_189_4 + _zz_when_ArraySlice_l173_189_8);
  assign _zz_when_ArraySlice_l173_189_4 = (_zz_when_ArraySlice_l173_189 - _zz_when_ArraySlice_l173_189_5);
  assign _zz_when_ArraySlice_l173_189_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_189_7);
  assign _zz_when_ArraySlice_l173_189_5 = {1'd0, _zz_when_ArraySlice_l173_189_6};
  assign _zz_when_ArraySlice_l173_189_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_189_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_190 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_190_1);
  assign _zz_when_ArraySlice_l165_190_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_190_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_190 = {1'd0, _zz_when_ArraySlice_l166_190_1};
  assign _zz_when_ArraySlice_l166_190_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_190_3);
  assign _zz_when_ArraySlice_l166_190_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_190_4);
  assign _zz_when_ArraySlice_l166_190_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_190 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_190 = (_zz_when_ArraySlice_l113_190_1 - _zz_when_ArraySlice_l113_190_4);
  assign _zz_when_ArraySlice_l113_190_1 = (_zz_when_ArraySlice_l113_190_2 + _zz_when_ArraySlice_l113_190_3);
  assign _zz_when_ArraySlice_l113_190_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_190_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_190_4 = {1'd0, _zz_when_ArraySlice_l112_190};
  assign _zz__zz_when_ArraySlice_l173_190 = (_zz__zz_when_ArraySlice_l173_190_1 + _zz__zz_when_ArraySlice_l173_190_2);
  assign _zz__zz_when_ArraySlice_l173_190_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_190_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_190_3 = {1'd0, _zz_when_ArraySlice_l112_190};
  assign _zz_when_ArraySlice_l118_190_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_190 = _zz_when_ArraySlice_l118_190_1[5:0];
  assign _zz_when_ArraySlice_l173_190_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_190_1 = {2'd0, _zz_when_ArraySlice_l173_190_2};
  assign _zz_when_ArraySlice_l173_190_3 = (_zz_when_ArraySlice_l173_190_4 + _zz_when_ArraySlice_l173_190_8);
  assign _zz_when_ArraySlice_l173_190_4 = (_zz_when_ArraySlice_l173_190 - _zz_when_ArraySlice_l173_190_5);
  assign _zz_when_ArraySlice_l173_190_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_190_7);
  assign _zz_when_ArraySlice_l173_190_5 = {1'd0, _zz_when_ArraySlice_l173_190_6};
  assign _zz_when_ArraySlice_l173_190_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_190_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_191 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_191_1);
  assign _zz_when_ArraySlice_l165_191_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_191_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_191 = {2'd0, _zz_when_ArraySlice_l166_191_1};
  assign _zz_when_ArraySlice_l166_191_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_191_3);
  assign _zz_when_ArraySlice_l166_191_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_191_4);
  assign _zz_when_ArraySlice_l166_191_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_191 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_191 = (_zz_when_ArraySlice_l113_191_1 - _zz_when_ArraySlice_l113_191_4);
  assign _zz_when_ArraySlice_l113_191_1 = (_zz_when_ArraySlice_l113_191_2 + _zz_when_ArraySlice_l113_191_3);
  assign _zz_when_ArraySlice_l113_191_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_191_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_191_4 = {1'd0, _zz_when_ArraySlice_l112_191};
  assign _zz__zz_when_ArraySlice_l173_191 = (_zz__zz_when_ArraySlice_l173_191_1 + _zz__zz_when_ArraySlice_l173_191_2);
  assign _zz__zz_when_ArraySlice_l173_191_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_191_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_191_3 = {1'd0, _zz_when_ArraySlice_l112_191};
  assign _zz_when_ArraySlice_l118_191_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_191 = _zz_when_ArraySlice_l118_191_1[5:0];
  assign _zz_when_ArraySlice_l173_191_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_191_1 = {3'd0, _zz_when_ArraySlice_l173_191_2};
  assign _zz_when_ArraySlice_l173_191_3 = (_zz_when_ArraySlice_l173_191_4 + _zz_when_ArraySlice_l173_191_8);
  assign _zz_when_ArraySlice_l173_191_4 = (_zz_when_ArraySlice_l173_191 - _zz_when_ArraySlice_l173_191_5);
  assign _zz_when_ArraySlice_l173_191_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_191_7);
  assign _zz_when_ArraySlice_l173_191_5 = {1'd0, _zz_when_ArraySlice_l173_191_6};
  assign _zz_when_ArraySlice_l173_191_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_191_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l421_7_1 = (_zz_when_ArraySlice_l421_7_2 + _zz_when_ArraySlice_l421_7_7);
  assign _zz_when_ArraySlice_l421_7_2 = (_zz_when_ArraySlice_l421_7_3 + _zz_when_ArraySlice_l421_7_5);
  assign _zz_when_ArraySlice_l421_7_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l421_7_4);
  assign _zz_when_ArraySlice_l421_7_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l421_7_6 = 1'b1;
  assign _zz_when_ArraySlice_l421_7_5 = {5'd0, _zz_when_ArraySlice_l421_7_6};
  assign _zz_when_ArraySlice_l421_7_7 = (bReg * 3'b111);
  assign _zz_selectReadFifo_7_25 = 1'b1;
  assign _zz_selectReadFifo_7_24 = {5'd0, _zz_selectReadFifo_7_25};
  assign _zz_when_ArraySlice_l425_7 = (_zz_when_ArraySlice_l425_7_1 % aReg);
  assign _zz_when_ArraySlice_l425_7_1 = (handshakeTimes_7_value + _zz_when_ArraySlice_l425_7_2);
  assign _zz_when_ArraySlice_l425_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l425_7_2 = {12'd0, _zz_when_ArraySlice_l425_7_3};
  assign _zz_when_ArraySlice_l436_7_1 = (_zz_when_ArraySlice_l436_7_2 - _zz_when_ArraySlice_l436_7_3);
  assign _zz_when_ArraySlice_l436_7 = {7'd0, _zz_when_ArraySlice_l436_7_1};
  assign _zz_when_ArraySlice_l436_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l436_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l436_7_3 = {5'd0, _zz_when_ArraySlice_l436_7_4};
  assign _zz__zz_when_ArraySlice_l94_23 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_23 = (_zz_when_ArraySlice_l95_23_1 - _zz_when_ArraySlice_l95_23_4);
  assign _zz_when_ArraySlice_l95_23_1 = (_zz_when_ArraySlice_l95_23_2 + _zz_when_ArraySlice_l95_23_3);
  assign _zz_when_ArraySlice_l95_23_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_23_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_23_4 = {1'd0, _zz_when_ArraySlice_l94_23};
  assign _zz__zz_when_ArraySlice_l437_7 = (_zz__zz_when_ArraySlice_l437_7_1 + _zz__zz_when_ArraySlice_l437_7_2);
  assign _zz__zz_when_ArraySlice_l437_7_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l437_7_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l437_7_3 = {1'd0, _zz_when_ArraySlice_l94_23};
  assign _zz_when_ArraySlice_l99_23_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_23 = _zz_when_ArraySlice_l99_23_1[5:0];
  assign _zz_when_ArraySlice_l437_7_1 = (outSliceNumb_7_value + _zz_when_ArraySlice_l437_7_2);
  assign _zz_when_ArraySlice_l437_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l437_7_2 = {6'd0, _zz_when_ArraySlice_l437_7_3};
  assign _zz_when_ArraySlice_l437_7_4 = (_zz_when_ArraySlice_l437_7 / aReg);
  assign _zz_selectReadFifo_7_26 = (selectReadFifo_7 - _zz_selectReadFifo_7_27);
  assign _zz_selectReadFifo_7_27 = {3'd0, bReg};
  assign _zz_selectReadFifo_7_29 = 1'b1;
  assign _zz_selectReadFifo_7_28 = {5'd0, _zz_selectReadFifo_7_29};
  assign _zz_when_ArraySlice_l165_192 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_192_1);
  assign _zz_when_ArraySlice_l165_192_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_192_1 = {3'd0, _zz_when_ArraySlice_l165_192_2};
  assign _zz_when_ArraySlice_l166_192 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_192_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_192_3);
  assign _zz_when_ArraySlice_l166_192_1 = {1'd0, _zz_when_ArraySlice_l166_192_2};
  assign _zz_when_ArraySlice_l166_192_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_192_4);
  assign _zz_when_ArraySlice_l166_192_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_192_4 = {3'd0, _zz_when_ArraySlice_l166_192_5};
  assign _zz__zz_when_ArraySlice_l112_192 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_192 = (_zz_when_ArraySlice_l113_192_1 - _zz_when_ArraySlice_l113_192_4);
  assign _zz_when_ArraySlice_l113_192_1 = (_zz_when_ArraySlice_l113_192_2 + _zz_when_ArraySlice_l113_192_3);
  assign _zz_when_ArraySlice_l113_192_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_192_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_192_4 = {1'd0, _zz_when_ArraySlice_l112_192};
  assign _zz__zz_when_ArraySlice_l173_192 = (_zz__zz_when_ArraySlice_l173_192_1 + _zz__zz_when_ArraySlice_l173_192_2);
  assign _zz__zz_when_ArraySlice_l173_192_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_192_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_192_3 = {1'd0, _zz_when_ArraySlice_l112_192};
  assign _zz_when_ArraySlice_l118_192_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_192 = _zz_when_ArraySlice_l118_192_1[5:0];
  assign _zz_when_ArraySlice_l173_192_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_192_2 = (_zz_when_ArraySlice_l173_192_3 + _zz_when_ArraySlice_l173_192_8);
  assign _zz_when_ArraySlice_l173_192_3 = (_zz_when_ArraySlice_l173_192 - _zz_when_ArraySlice_l173_192_4);
  assign _zz_when_ArraySlice_l173_192_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_192_6);
  assign _zz_when_ArraySlice_l173_192_4 = {1'd0, _zz_when_ArraySlice_l173_192_5};
  assign _zz_when_ArraySlice_l173_192_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_192_6 = {3'd0, _zz_when_ArraySlice_l173_192_7};
  assign _zz_when_ArraySlice_l173_192_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_193 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_193_1);
  assign _zz_when_ArraySlice_l165_193_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_193_1 = {2'd0, _zz_when_ArraySlice_l165_193_2};
  assign _zz_when_ArraySlice_l166_193 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_193_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_193_2);
  assign _zz_when_ArraySlice_l166_193_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_193_3);
  assign _zz_when_ArraySlice_l166_193_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_193_3 = {2'd0, _zz_when_ArraySlice_l166_193_4};
  assign _zz__zz_when_ArraySlice_l112_193 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_193 = (_zz_when_ArraySlice_l113_193_1 - _zz_when_ArraySlice_l113_193_4);
  assign _zz_when_ArraySlice_l113_193_1 = (_zz_when_ArraySlice_l113_193_2 + _zz_when_ArraySlice_l113_193_3);
  assign _zz_when_ArraySlice_l113_193_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_193_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_193_4 = {1'd0, _zz_when_ArraySlice_l112_193};
  assign _zz__zz_when_ArraySlice_l173_193 = (_zz__zz_when_ArraySlice_l173_193_1 + _zz__zz_when_ArraySlice_l173_193_2);
  assign _zz__zz_when_ArraySlice_l173_193_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_193_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_193_3 = {1'd0, _zz_when_ArraySlice_l112_193};
  assign _zz_when_ArraySlice_l118_193_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_193 = _zz_when_ArraySlice_l118_193_1[5:0];
  assign _zz_when_ArraySlice_l173_193_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_193_1 = {1'd0, _zz_when_ArraySlice_l173_193_2};
  assign _zz_when_ArraySlice_l173_193_3 = (_zz_when_ArraySlice_l173_193_4 + _zz_when_ArraySlice_l173_193_9);
  assign _zz_when_ArraySlice_l173_193_4 = (_zz_when_ArraySlice_l173_193 - _zz_when_ArraySlice_l173_193_5);
  assign _zz_when_ArraySlice_l173_193_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_193_7);
  assign _zz_when_ArraySlice_l173_193_5 = {1'd0, _zz_when_ArraySlice_l173_193_6};
  assign _zz_when_ArraySlice_l173_193_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_193_7 = {2'd0, _zz_when_ArraySlice_l173_193_8};
  assign _zz_when_ArraySlice_l173_193_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_194 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_194_1);
  assign _zz_when_ArraySlice_l165_194_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_194_1 = {1'd0, _zz_when_ArraySlice_l165_194_2};
  assign _zz_when_ArraySlice_l166_194 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_194_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_194_2);
  assign _zz_when_ArraySlice_l166_194_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_194_3);
  assign _zz_when_ArraySlice_l166_194_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_194_3 = {1'd0, _zz_when_ArraySlice_l166_194_4};
  assign _zz__zz_when_ArraySlice_l112_194 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_194 = (_zz_when_ArraySlice_l113_194_1 - _zz_when_ArraySlice_l113_194_4);
  assign _zz_when_ArraySlice_l113_194_1 = (_zz_when_ArraySlice_l113_194_2 + _zz_when_ArraySlice_l113_194_3);
  assign _zz_when_ArraySlice_l113_194_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_194_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_194_4 = {1'd0, _zz_when_ArraySlice_l112_194};
  assign _zz__zz_when_ArraySlice_l173_194 = (_zz__zz_when_ArraySlice_l173_194_1 + _zz__zz_when_ArraySlice_l173_194_2);
  assign _zz__zz_when_ArraySlice_l173_194_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_194_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_194_3 = {1'd0, _zz_when_ArraySlice_l112_194};
  assign _zz_when_ArraySlice_l118_194_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_194 = _zz_when_ArraySlice_l118_194_1[5:0];
  assign _zz_when_ArraySlice_l173_194_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_194_1 = {1'd0, _zz_when_ArraySlice_l173_194_2};
  assign _zz_when_ArraySlice_l173_194_3 = (_zz_when_ArraySlice_l173_194_4 + _zz_when_ArraySlice_l173_194_9);
  assign _zz_when_ArraySlice_l173_194_4 = (_zz_when_ArraySlice_l173_194 - _zz_when_ArraySlice_l173_194_5);
  assign _zz_when_ArraySlice_l173_194_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_194_7);
  assign _zz_when_ArraySlice_l173_194_5 = {1'd0, _zz_when_ArraySlice_l173_194_6};
  assign _zz_when_ArraySlice_l173_194_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_194_7 = {1'd0, _zz_when_ArraySlice_l173_194_8};
  assign _zz_when_ArraySlice_l173_194_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_195 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_195_1);
  assign _zz_when_ArraySlice_l165_195_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_195_1 = {1'd0, _zz_when_ArraySlice_l165_195_2};
  assign _zz_when_ArraySlice_l166_195 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_195_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_195_2);
  assign _zz_when_ArraySlice_l166_195_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_195_3);
  assign _zz_when_ArraySlice_l166_195_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_195_3 = {1'd0, _zz_when_ArraySlice_l166_195_4};
  assign _zz__zz_when_ArraySlice_l112_195 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_195 = (_zz_when_ArraySlice_l113_195_1 - _zz_when_ArraySlice_l113_195_4);
  assign _zz_when_ArraySlice_l113_195_1 = (_zz_when_ArraySlice_l113_195_2 + _zz_when_ArraySlice_l113_195_3);
  assign _zz_when_ArraySlice_l113_195_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_195_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_195_4 = {1'd0, _zz_when_ArraySlice_l112_195};
  assign _zz__zz_when_ArraySlice_l173_195 = (_zz__zz_when_ArraySlice_l173_195_1 + _zz__zz_when_ArraySlice_l173_195_2);
  assign _zz__zz_when_ArraySlice_l173_195_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_195_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_195_3 = {1'd0, _zz_when_ArraySlice_l112_195};
  assign _zz_when_ArraySlice_l118_195_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_195 = _zz_when_ArraySlice_l118_195_1[5:0];
  assign _zz_when_ArraySlice_l173_195_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_195_1 = {1'd0, _zz_when_ArraySlice_l173_195_2};
  assign _zz_when_ArraySlice_l173_195_3 = (_zz_when_ArraySlice_l173_195_4 + _zz_when_ArraySlice_l173_195_9);
  assign _zz_when_ArraySlice_l173_195_4 = (_zz_when_ArraySlice_l173_195 - _zz_when_ArraySlice_l173_195_5);
  assign _zz_when_ArraySlice_l173_195_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_195_7);
  assign _zz_when_ArraySlice_l173_195_5 = {1'd0, _zz_when_ArraySlice_l173_195_6};
  assign _zz_when_ArraySlice_l173_195_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_195_7 = {1'd0, _zz_when_ArraySlice_l173_195_8};
  assign _zz_when_ArraySlice_l173_195_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_196 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_196_1);
  assign _zz_when_ArraySlice_l165_196_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_196 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_196_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_196_2);
  assign _zz_when_ArraySlice_l166_196_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_196_3);
  assign _zz_when_ArraySlice_l166_196_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_196 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_196 = (_zz_when_ArraySlice_l113_196_1 - _zz_when_ArraySlice_l113_196_4);
  assign _zz_when_ArraySlice_l113_196_1 = (_zz_when_ArraySlice_l113_196_2 + _zz_when_ArraySlice_l113_196_3);
  assign _zz_when_ArraySlice_l113_196_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_196_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_196_4 = {1'd0, _zz_when_ArraySlice_l112_196};
  assign _zz__zz_when_ArraySlice_l173_196 = (_zz__zz_when_ArraySlice_l173_196_1 + _zz__zz_when_ArraySlice_l173_196_2);
  assign _zz__zz_when_ArraySlice_l173_196_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_196_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_196_3 = {1'd0, _zz_when_ArraySlice_l112_196};
  assign _zz_when_ArraySlice_l118_196_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_196 = _zz_when_ArraySlice_l118_196_1[5:0];
  assign _zz_when_ArraySlice_l173_196_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_196_1 = {1'd0, _zz_when_ArraySlice_l173_196_2};
  assign _zz_when_ArraySlice_l173_196_3 = (_zz_when_ArraySlice_l173_196_4 + _zz_when_ArraySlice_l173_196_8);
  assign _zz_when_ArraySlice_l173_196_4 = (_zz_when_ArraySlice_l173_196 - _zz_when_ArraySlice_l173_196_5);
  assign _zz_when_ArraySlice_l173_196_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_196_7);
  assign _zz_when_ArraySlice_l173_196_5 = {1'd0, _zz_when_ArraySlice_l173_196_6};
  assign _zz_when_ArraySlice_l173_196_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_196_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_197 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_197_1);
  assign _zz_when_ArraySlice_l165_197_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_197_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_197 = {1'd0, _zz_when_ArraySlice_l166_197_1};
  assign _zz_when_ArraySlice_l166_197_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_197_3);
  assign _zz_when_ArraySlice_l166_197_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_197_4);
  assign _zz_when_ArraySlice_l166_197_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_197 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_197 = (_zz_when_ArraySlice_l113_197_1 - _zz_when_ArraySlice_l113_197_4);
  assign _zz_when_ArraySlice_l113_197_1 = (_zz_when_ArraySlice_l113_197_2 + _zz_when_ArraySlice_l113_197_3);
  assign _zz_when_ArraySlice_l113_197_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_197_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_197_4 = {1'd0, _zz_when_ArraySlice_l112_197};
  assign _zz__zz_when_ArraySlice_l173_197 = (_zz__zz_when_ArraySlice_l173_197_1 + _zz__zz_when_ArraySlice_l173_197_2);
  assign _zz__zz_when_ArraySlice_l173_197_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_197_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_197_3 = {1'd0, _zz_when_ArraySlice_l112_197};
  assign _zz_when_ArraySlice_l118_197_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_197 = _zz_when_ArraySlice_l118_197_1[5:0];
  assign _zz_when_ArraySlice_l173_197_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_197_1 = {2'd0, _zz_when_ArraySlice_l173_197_2};
  assign _zz_when_ArraySlice_l173_197_3 = (_zz_when_ArraySlice_l173_197_4 + _zz_when_ArraySlice_l173_197_8);
  assign _zz_when_ArraySlice_l173_197_4 = (_zz_when_ArraySlice_l173_197 - _zz_when_ArraySlice_l173_197_5);
  assign _zz_when_ArraySlice_l173_197_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_197_7);
  assign _zz_when_ArraySlice_l173_197_5 = {1'd0, _zz_when_ArraySlice_l173_197_6};
  assign _zz_when_ArraySlice_l173_197_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_197_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_198 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_198_1);
  assign _zz_when_ArraySlice_l165_198_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_198_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_198 = {1'd0, _zz_when_ArraySlice_l166_198_1};
  assign _zz_when_ArraySlice_l166_198_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_198_3);
  assign _zz_when_ArraySlice_l166_198_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_198_4);
  assign _zz_when_ArraySlice_l166_198_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_198 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_198 = (_zz_when_ArraySlice_l113_198_1 - _zz_when_ArraySlice_l113_198_4);
  assign _zz_when_ArraySlice_l113_198_1 = (_zz_when_ArraySlice_l113_198_2 + _zz_when_ArraySlice_l113_198_3);
  assign _zz_when_ArraySlice_l113_198_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_198_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_198_4 = {1'd0, _zz_when_ArraySlice_l112_198};
  assign _zz__zz_when_ArraySlice_l173_198 = (_zz__zz_when_ArraySlice_l173_198_1 + _zz__zz_when_ArraySlice_l173_198_2);
  assign _zz__zz_when_ArraySlice_l173_198_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_198_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_198_3 = {1'd0, _zz_when_ArraySlice_l112_198};
  assign _zz_when_ArraySlice_l118_198_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_198 = _zz_when_ArraySlice_l118_198_1[5:0];
  assign _zz_when_ArraySlice_l173_198_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_198_1 = {2'd0, _zz_when_ArraySlice_l173_198_2};
  assign _zz_when_ArraySlice_l173_198_3 = (_zz_when_ArraySlice_l173_198_4 + _zz_when_ArraySlice_l173_198_8);
  assign _zz_when_ArraySlice_l173_198_4 = (_zz_when_ArraySlice_l173_198 - _zz_when_ArraySlice_l173_198_5);
  assign _zz_when_ArraySlice_l173_198_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_198_7);
  assign _zz_when_ArraySlice_l173_198_5 = {1'd0, _zz_when_ArraySlice_l173_198_6};
  assign _zz_when_ArraySlice_l173_198_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_198_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_199 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_199_1);
  assign _zz_when_ArraySlice_l165_199_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_199_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_199 = {2'd0, _zz_when_ArraySlice_l166_199_1};
  assign _zz_when_ArraySlice_l166_199_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_199_3);
  assign _zz_when_ArraySlice_l166_199_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_199_4);
  assign _zz_when_ArraySlice_l166_199_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_199 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_199 = (_zz_when_ArraySlice_l113_199_1 - _zz_when_ArraySlice_l113_199_4);
  assign _zz_when_ArraySlice_l113_199_1 = (_zz_when_ArraySlice_l113_199_2 + _zz_when_ArraySlice_l113_199_3);
  assign _zz_when_ArraySlice_l113_199_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_199_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_199_4 = {1'd0, _zz_when_ArraySlice_l112_199};
  assign _zz__zz_when_ArraySlice_l173_199 = (_zz__zz_when_ArraySlice_l173_199_1 + _zz__zz_when_ArraySlice_l173_199_2);
  assign _zz__zz_when_ArraySlice_l173_199_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_199_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_199_3 = {1'd0, _zz_when_ArraySlice_l112_199};
  assign _zz_when_ArraySlice_l118_199_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_199 = _zz_when_ArraySlice_l118_199_1[5:0];
  assign _zz_when_ArraySlice_l173_199_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_199_1 = {3'd0, _zz_when_ArraySlice_l173_199_2};
  assign _zz_when_ArraySlice_l173_199_3 = (_zz_when_ArraySlice_l173_199_4 + _zz_when_ArraySlice_l173_199_8);
  assign _zz_when_ArraySlice_l173_199_4 = (_zz_when_ArraySlice_l173_199 - _zz_when_ArraySlice_l173_199_5);
  assign _zz_when_ArraySlice_l173_199_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_199_7);
  assign _zz_when_ArraySlice_l173_199_5 = {1'd0, _zz_when_ArraySlice_l173_199_6};
  assign _zz_when_ArraySlice_l173_199_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_199_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_7_31 = 1'b1;
  assign _zz_selectReadFifo_7_30 = {5'd0, _zz_selectReadFifo_7_31};
  assign _zz_when_ArraySlice_l448_7 = (_zz_when_ArraySlice_l448_7_1 % aReg);
  assign _zz_when_ArraySlice_l448_7_1 = (handshakeTimes_7_value + _zz_when_ArraySlice_l448_7_2);
  assign _zz_when_ArraySlice_l448_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l448_7_2 = {12'd0, _zz_when_ArraySlice_l448_7_3};
  assign _zz_when_ArraySlice_l434_7 = (selectReadFifo_7 + _zz_when_ArraySlice_l434_7_1);
  assign _zz_when_ArraySlice_l434_7_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l455_7_1 = (_zz_when_ArraySlice_l455_7_2 - _zz_when_ArraySlice_l455_7_3);
  assign _zz_when_ArraySlice_l455_7 = {7'd0, _zz_when_ArraySlice_l455_7_1};
  assign _zz_when_ArraySlice_l455_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l455_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l455_7_3 = {5'd0, _zz_when_ArraySlice_l455_7_4};
  assign _zz_when_ArraySlice_l165_200 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_200_1);
  assign _zz_when_ArraySlice_l165_200_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_200_1 = {3'd0, _zz_when_ArraySlice_l165_200_2};
  assign _zz_when_ArraySlice_l166_200 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_200_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_200_3);
  assign _zz_when_ArraySlice_l166_200_1 = {1'd0, _zz_when_ArraySlice_l166_200_2};
  assign _zz_when_ArraySlice_l166_200_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_200_4);
  assign _zz_when_ArraySlice_l166_200_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_200_4 = {3'd0, _zz_when_ArraySlice_l166_200_5};
  assign _zz__zz_when_ArraySlice_l112_200 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_200 = (_zz_when_ArraySlice_l113_200_1 - _zz_when_ArraySlice_l113_200_4);
  assign _zz_when_ArraySlice_l113_200_1 = (_zz_when_ArraySlice_l113_200_2 + _zz_when_ArraySlice_l113_200_3);
  assign _zz_when_ArraySlice_l113_200_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_200_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_200_4 = {1'd0, _zz_when_ArraySlice_l112_200};
  assign _zz__zz_when_ArraySlice_l173_200 = (_zz__zz_when_ArraySlice_l173_200_1 + _zz__zz_when_ArraySlice_l173_200_2);
  assign _zz__zz_when_ArraySlice_l173_200_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_200_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_200_3 = {1'd0, _zz_when_ArraySlice_l112_200};
  assign _zz_when_ArraySlice_l118_200_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_200 = _zz_when_ArraySlice_l118_200_1[5:0];
  assign _zz_when_ArraySlice_l173_200_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_200_2 = (_zz_when_ArraySlice_l173_200_3 + _zz_when_ArraySlice_l173_200_8);
  assign _zz_when_ArraySlice_l173_200_3 = (_zz_when_ArraySlice_l173_200 - _zz_when_ArraySlice_l173_200_4);
  assign _zz_when_ArraySlice_l173_200_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_200_6);
  assign _zz_when_ArraySlice_l173_200_4 = {1'd0, _zz_when_ArraySlice_l173_200_5};
  assign _zz_when_ArraySlice_l173_200_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_200_6 = {3'd0, _zz_when_ArraySlice_l173_200_7};
  assign _zz_when_ArraySlice_l173_200_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_201 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_201_1);
  assign _zz_when_ArraySlice_l165_201_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_201_1 = {2'd0, _zz_when_ArraySlice_l165_201_2};
  assign _zz_when_ArraySlice_l166_201 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_201_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_201_2);
  assign _zz_when_ArraySlice_l166_201_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_201_3);
  assign _zz_when_ArraySlice_l166_201_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_201_3 = {2'd0, _zz_when_ArraySlice_l166_201_4};
  assign _zz__zz_when_ArraySlice_l112_201 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_201 = (_zz_when_ArraySlice_l113_201_1 - _zz_when_ArraySlice_l113_201_4);
  assign _zz_when_ArraySlice_l113_201_1 = (_zz_when_ArraySlice_l113_201_2 + _zz_when_ArraySlice_l113_201_3);
  assign _zz_when_ArraySlice_l113_201_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_201_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_201_4 = {1'd0, _zz_when_ArraySlice_l112_201};
  assign _zz__zz_when_ArraySlice_l173_201 = (_zz__zz_when_ArraySlice_l173_201_1 + _zz__zz_when_ArraySlice_l173_201_2);
  assign _zz__zz_when_ArraySlice_l173_201_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_201_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_201_3 = {1'd0, _zz_when_ArraySlice_l112_201};
  assign _zz_when_ArraySlice_l118_201_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_201 = _zz_when_ArraySlice_l118_201_1[5:0];
  assign _zz_when_ArraySlice_l173_201_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_201_1 = {1'd0, _zz_when_ArraySlice_l173_201_2};
  assign _zz_when_ArraySlice_l173_201_3 = (_zz_when_ArraySlice_l173_201_4 + _zz_when_ArraySlice_l173_201_9);
  assign _zz_when_ArraySlice_l173_201_4 = (_zz_when_ArraySlice_l173_201 - _zz_when_ArraySlice_l173_201_5);
  assign _zz_when_ArraySlice_l173_201_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_201_7);
  assign _zz_when_ArraySlice_l173_201_5 = {1'd0, _zz_when_ArraySlice_l173_201_6};
  assign _zz_when_ArraySlice_l173_201_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_201_7 = {2'd0, _zz_when_ArraySlice_l173_201_8};
  assign _zz_when_ArraySlice_l173_201_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_202 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_202_1);
  assign _zz_when_ArraySlice_l165_202_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_202_1 = {1'd0, _zz_when_ArraySlice_l165_202_2};
  assign _zz_when_ArraySlice_l166_202 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_202_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_202_2);
  assign _zz_when_ArraySlice_l166_202_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_202_3);
  assign _zz_when_ArraySlice_l166_202_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_202_3 = {1'd0, _zz_when_ArraySlice_l166_202_4};
  assign _zz__zz_when_ArraySlice_l112_202 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_202 = (_zz_when_ArraySlice_l113_202_1 - _zz_when_ArraySlice_l113_202_4);
  assign _zz_when_ArraySlice_l113_202_1 = (_zz_when_ArraySlice_l113_202_2 + _zz_when_ArraySlice_l113_202_3);
  assign _zz_when_ArraySlice_l113_202_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_202_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_202_4 = {1'd0, _zz_when_ArraySlice_l112_202};
  assign _zz__zz_when_ArraySlice_l173_202 = (_zz__zz_when_ArraySlice_l173_202_1 + _zz__zz_when_ArraySlice_l173_202_2);
  assign _zz__zz_when_ArraySlice_l173_202_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_202_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_202_3 = {1'd0, _zz_when_ArraySlice_l112_202};
  assign _zz_when_ArraySlice_l118_202_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_202 = _zz_when_ArraySlice_l118_202_1[5:0];
  assign _zz_when_ArraySlice_l173_202_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_202_1 = {1'd0, _zz_when_ArraySlice_l173_202_2};
  assign _zz_when_ArraySlice_l173_202_3 = (_zz_when_ArraySlice_l173_202_4 + _zz_when_ArraySlice_l173_202_9);
  assign _zz_when_ArraySlice_l173_202_4 = (_zz_when_ArraySlice_l173_202 - _zz_when_ArraySlice_l173_202_5);
  assign _zz_when_ArraySlice_l173_202_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_202_7);
  assign _zz_when_ArraySlice_l173_202_5 = {1'd0, _zz_when_ArraySlice_l173_202_6};
  assign _zz_when_ArraySlice_l173_202_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_202_7 = {1'd0, _zz_when_ArraySlice_l173_202_8};
  assign _zz_when_ArraySlice_l173_202_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_203 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_203_1);
  assign _zz_when_ArraySlice_l165_203_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_203_1 = {1'd0, _zz_when_ArraySlice_l165_203_2};
  assign _zz_when_ArraySlice_l166_203 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_203_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_203_2);
  assign _zz_when_ArraySlice_l166_203_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_203_3);
  assign _zz_when_ArraySlice_l166_203_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_203_3 = {1'd0, _zz_when_ArraySlice_l166_203_4};
  assign _zz__zz_when_ArraySlice_l112_203 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_203 = (_zz_when_ArraySlice_l113_203_1 - _zz_when_ArraySlice_l113_203_4);
  assign _zz_when_ArraySlice_l113_203_1 = (_zz_when_ArraySlice_l113_203_2 + _zz_when_ArraySlice_l113_203_3);
  assign _zz_when_ArraySlice_l113_203_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_203_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_203_4 = {1'd0, _zz_when_ArraySlice_l112_203};
  assign _zz__zz_when_ArraySlice_l173_203 = (_zz__zz_when_ArraySlice_l173_203_1 + _zz__zz_when_ArraySlice_l173_203_2);
  assign _zz__zz_when_ArraySlice_l173_203_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_203_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_203_3 = {1'd0, _zz_when_ArraySlice_l112_203};
  assign _zz_when_ArraySlice_l118_203_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_203 = _zz_when_ArraySlice_l118_203_1[5:0];
  assign _zz_when_ArraySlice_l173_203_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_203_1 = {1'd0, _zz_when_ArraySlice_l173_203_2};
  assign _zz_when_ArraySlice_l173_203_3 = (_zz_when_ArraySlice_l173_203_4 + _zz_when_ArraySlice_l173_203_9);
  assign _zz_when_ArraySlice_l173_203_4 = (_zz_when_ArraySlice_l173_203 - _zz_when_ArraySlice_l173_203_5);
  assign _zz_when_ArraySlice_l173_203_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_203_7);
  assign _zz_when_ArraySlice_l173_203_5 = {1'd0, _zz_when_ArraySlice_l173_203_6};
  assign _zz_when_ArraySlice_l173_203_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_203_7 = {1'd0, _zz_when_ArraySlice_l173_203_8};
  assign _zz_when_ArraySlice_l173_203_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_204 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_204_1);
  assign _zz_when_ArraySlice_l165_204_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_204 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_204_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_204_2);
  assign _zz_when_ArraySlice_l166_204_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_204_3);
  assign _zz_when_ArraySlice_l166_204_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_204 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_204 = (_zz_when_ArraySlice_l113_204_1 - _zz_when_ArraySlice_l113_204_4);
  assign _zz_when_ArraySlice_l113_204_1 = (_zz_when_ArraySlice_l113_204_2 + _zz_when_ArraySlice_l113_204_3);
  assign _zz_when_ArraySlice_l113_204_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_204_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_204_4 = {1'd0, _zz_when_ArraySlice_l112_204};
  assign _zz__zz_when_ArraySlice_l173_204 = (_zz__zz_when_ArraySlice_l173_204_1 + _zz__zz_when_ArraySlice_l173_204_2);
  assign _zz__zz_when_ArraySlice_l173_204_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_204_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_204_3 = {1'd0, _zz_when_ArraySlice_l112_204};
  assign _zz_when_ArraySlice_l118_204_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_204 = _zz_when_ArraySlice_l118_204_1[5:0];
  assign _zz_when_ArraySlice_l173_204_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_204_1 = {1'd0, _zz_when_ArraySlice_l173_204_2};
  assign _zz_when_ArraySlice_l173_204_3 = (_zz_when_ArraySlice_l173_204_4 + _zz_when_ArraySlice_l173_204_8);
  assign _zz_when_ArraySlice_l173_204_4 = (_zz_when_ArraySlice_l173_204 - _zz_when_ArraySlice_l173_204_5);
  assign _zz_when_ArraySlice_l173_204_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_204_7);
  assign _zz_when_ArraySlice_l173_204_5 = {1'd0, _zz_when_ArraySlice_l173_204_6};
  assign _zz_when_ArraySlice_l173_204_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_204_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_205 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_205_1);
  assign _zz_when_ArraySlice_l165_205_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_205_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_205 = {1'd0, _zz_when_ArraySlice_l166_205_1};
  assign _zz_when_ArraySlice_l166_205_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_205_3);
  assign _zz_when_ArraySlice_l166_205_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_205_4);
  assign _zz_when_ArraySlice_l166_205_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_205 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_205 = (_zz_when_ArraySlice_l113_205_1 - _zz_when_ArraySlice_l113_205_4);
  assign _zz_when_ArraySlice_l113_205_1 = (_zz_when_ArraySlice_l113_205_2 + _zz_when_ArraySlice_l113_205_3);
  assign _zz_when_ArraySlice_l113_205_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_205_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_205_4 = {1'd0, _zz_when_ArraySlice_l112_205};
  assign _zz__zz_when_ArraySlice_l173_205 = (_zz__zz_when_ArraySlice_l173_205_1 + _zz__zz_when_ArraySlice_l173_205_2);
  assign _zz__zz_when_ArraySlice_l173_205_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_205_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_205_3 = {1'd0, _zz_when_ArraySlice_l112_205};
  assign _zz_when_ArraySlice_l118_205_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_205 = _zz_when_ArraySlice_l118_205_1[5:0];
  assign _zz_when_ArraySlice_l173_205_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_205_1 = {2'd0, _zz_when_ArraySlice_l173_205_2};
  assign _zz_when_ArraySlice_l173_205_3 = (_zz_when_ArraySlice_l173_205_4 + _zz_when_ArraySlice_l173_205_8);
  assign _zz_when_ArraySlice_l173_205_4 = (_zz_when_ArraySlice_l173_205 - _zz_when_ArraySlice_l173_205_5);
  assign _zz_when_ArraySlice_l173_205_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_205_7);
  assign _zz_when_ArraySlice_l173_205_5 = {1'd0, _zz_when_ArraySlice_l173_205_6};
  assign _zz_when_ArraySlice_l173_205_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_205_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_206 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_206_1);
  assign _zz_when_ArraySlice_l165_206_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_206_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_206 = {1'd0, _zz_when_ArraySlice_l166_206_1};
  assign _zz_when_ArraySlice_l166_206_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_206_3);
  assign _zz_when_ArraySlice_l166_206_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_206_4);
  assign _zz_when_ArraySlice_l166_206_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_206 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_206 = (_zz_when_ArraySlice_l113_206_1 - _zz_when_ArraySlice_l113_206_4);
  assign _zz_when_ArraySlice_l113_206_1 = (_zz_when_ArraySlice_l113_206_2 + _zz_when_ArraySlice_l113_206_3);
  assign _zz_when_ArraySlice_l113_206_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_206_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_206_4 = {1'd0, _zz_when_ArraySlice_l112_206};
  assign _zz__zz_when_ArraySlice_l173_206 = (_zz__zz_when_ArraySlice_l173_206_1 + _zz__zz_when_ArraySlice_l173_206_2);
  assign _zz__zz_when_ArraySlice_l173_206_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_206_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_206_3 = {1'd0, _zz_when_ArraySlice_l112_206};
  assign _zz_when_ArraySlice_l118_206_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_206 = _zz_when_ArraySlice_l118_206_1[5:0];
  assign _zz_when_ArraySlice_l173_206_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_206_1 = {2'd0, _zz_when_ArraySlice_l173_206_2};
  assign _zz_when_ArraySlice_l173_206_3 = (_zz_when_ArraySlice_l173_206_4 + _zz_when_ArraySlice_l173_206_8);
  assign _zz_when_ArraySlice_l173_206_4 = (_zz_when_ArraySlice_l173_206 - _zz_when_ArraySlice_l173_206_5);
  assign _zz_when_ArraySlice_l173_206_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_206_7);
  assign _zz_when_ArraySlice_l173_206_5 = {1'd0, _zz_when_ArraySlice_l173_206_6};
  assign _zz_when_ArraySlice_l173_206_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_206_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_207 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_207_1);
  assign _zz_when_ArraySlice_l165_207_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_207_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_207 = {2'd0, _zz_when_ArraySlice_l166_207_1};
  assign _zz_when_ArraySlice_l166_207_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_207_3);
  assign _zz_when_ArraySlice_l166_207_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_207_4);
  assign _zz_when_ArraySlice_l166_207_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_207 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_207 = (_zz_when_ArraySlice_l113_207_1 - _zz_when_ArraySlice_l113_207_4);
  assign _zz_when_ArraySlice_l113_207_1 = (_zz_when_ArraySlice_l113_207_2 + _zz_when_ArraySlice_l113_207_3);
  assign _zz_when_ArraySlice_l113_207_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_207_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_207_4 = {1'd0, _zz_when_ArraySlice_l112_207};
  assign _zz__zz_when_ArraySlice_l173_207 = (_zz__zz_when_ArraySlice_l173_207_1 + _zz__zz_when_ArraySlice_l173_207_2);
  assign _zz__zz_when_ArraySlice_l173_207_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_207_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_207_3 = {1'd0, _zz_when_ArraySlice_l112_207};
  assign _zz_when_ArraySlice_l118_207_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_207 = _zz_when_ArraySlice_l118_207_1[5:0];
  assign _zz_when_ArraySlice_l173_207_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_207_1 = {3'd0, _zz_when_ArraySlice_l173_207_2};
  assign _zz_when_ArraySlice_l173_207_3 = (_zz_when_ArraySlice_l173_207_4 + _zz_when_ArraySlice_l173_207_8);
  assign _zz_when_ArraySlice_l173_207_4 = (_zz_when_ArraySlice_l173_207 - _zz_when_ArraySlice_l173_207_5);
  assign _zz_when_ArraySlice_l173_207_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_207_7);
  assign _zz_when_ArraySlice_l173_207_5 = {1'd0, _zz_when_ArraySlice_l173_207_6};
  assign _zz_when_ArraySlice_l173_207_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_207_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l240 = (selectReadFifo_0 + _zz_when_ArraySlice_l240_1);
  assign _zz_when_ArraySlice_l240_2 = 3'b000;
  assign _zz_when_ArraySlice_l240_1 = {3'd0, _zz_when_ArraySlice_l240_2};
  assign _zz_when_ArraySlice_l241_1 = (selectReadFifo_0 + _zz_when_ArraySlice_l241_2);
  assign _zz_when_ArraySlice_l241_3 = 3'b000;
  assign _zz_when_ArraySlice_l241_2 = {3'd0, _zz_when_ArraySlice_l241_3};
  assign _zz__zz_outputStreamArrayData_0_valid_1_2 = 3'b000;
  assign _zz__zz_outputStreamArrayData_0_valid_1_1 = {3'd0, _zz__zz_outputStreamArrayData_0_valid_1_2};
  assign _zz_when_ArraySlice_l247_1 = 1'b1;
  assign _zz_when_ArraySlice_l247 = {6'd0, _zz_when_ArraySlice_l247_1};
  assign _zz_when_ArraySlice_l247_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l247_4);
  assign _zz_when_ArraySlice_l247_5 = 3'b000;
  assign _zz_when_ArraySlice_l247_4 = {3'd0, _zz_when_ArraySlice_l247_5};
  assign _zz_when_ArraySlice_l248_1 = (_zz_when_ArraySlice_l248_2 - _zz_when_ArraySlice_l248_3);
  assign _zz_when_ArraySlice_l248 = {7'd0, _zz_when_ArraySlice_l248_1};
  assign _zz_when_ArraySlice_l248_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l248_4 = 1'b1;
  assign _zz_when_ArraySlice_l248_3 = {5'd0, _zz_when_ArraySlice_l248_4};
  assign _zz_selectReadFifo_0_32 = (selectReadFifo_0 - _zz_selectReadFifo_0_33);
  assign _zz_selectReadFifo_0_33 = {3'd0, bReg};
  assign _zz_selectReadFifo_0_35 = 1'b1;
  assign _zz_selectReadFifo_0_34 = {5'd0, _zz_selectReadFifo_0_35};
  assign _zz_selectReadFifo_0_37 = 1'b1;
  assign _zz_selectReadFifo_0_36 = {5'd0, _zz_selectReadFifo_0_37};
  assign _zz_when_ArraySlice_l251 = (_zz_when_ArraySlice_l251_1 % aReg);
  assign _zz_when_ArraySlice_l251_1 = (handshakeTimes_0_value + _zz_when_ArraySlice_l251_2);
  assign _zz_when_ArraySlice_l251_3 = 1'b1;
  assign _zz_when_ArraySlice_l251_2 = {12'd0, _zz_when_ArraySlice_l251_3};
  assign _zz_when_ArraySlice_l256_1 = (selectReadFifo_0 + _zz_when_ArraySlice_l256_2);
  assign _zz_when_ArraySlice_l256_3 = 3'b000;
  assign _zz_when_ArraySlice_l256_2 = {3'd0, _zz_when_ArraySlice_l256_3};
  assign _zz_when_ArraySlice_l256_5 = 1'b1;
  assign _zz_when_ArraySlice_l256_4 = {6'd0, _zz_when_ArraySlice_l256_5};
  assign _zz_when_ArraySlice_l257_1 = (_zz_when_ArraySlice_l257_2 - _zz_when_ArraySlice_l257_3);
  assign _zz_when_ArraySlice_l257 = {7'd0, _zz_when_ArraySlice_l257_1};
  assign _zz_when_ArraySlice_l257_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l257_4 = 1'b1;
  assign _zz_when_ArraySlice_l257_3 = {5'd0, _zz_when_ArraySlice_l257_4};
  assign _zz__zz_when_ArraySlice_l94_24 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_24 = (_zz_when_ArraySlice_l95_24_1 - _zz_when_ArraySlice_l95_24_4);
  assign _zz_when_ArraySlice_l95_24_1 = (_zz_when_ArraySlice_l95_24_2 + _zz_when_ArraySlice_l95_24_3);
  assign _zz_when_ArraySlice_l95_24_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_24_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_24_4 = {1'd0, _zz_when_ArraySlice_l94_24};
  assign _zz__zz_when_ArraySlice_l259 = (_zz__zz_when_ArraySlice_l259_1 + _zz__zz_when_ArraySlice_l259_2);
  assign _zz__zz_when_ArraySlice_l259_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l259_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l259_3 = {1'd0, _zz_when_ArraySlice_l94_24};
  assign _zz_when_ArraySlice_l99_24_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_24 = _zz_when_ArraySlice_l99_24_1[5:0];
  assign _zz_when_ArraySlice_l259_8 = (outSliceNumb_0_value + _zz_when_ArraySlice_l259_9);
  assign _zz_when_ArraySlice_l259_10 = 1'b1;
  assign _zz_when_ArraySlice_l259_9 = {6'd0, _zz_when_ArraySlice_l259_10};
  assign _zz_when_ArraySlice_l259_11 = (_zz_when_ArraySlice_l259 / aReg);
  assign _zz_selectReadFifo_0_38 = (selectReadFifo_0 - _zz_selectReadFifo_0_39);
  assign _zz_selectReadFifo_0_39 = {3'd0, bReg};
  assign _zz_selectReadFifo_0_41 = 1'b1;
  assign _zz_selectReadFifo_0_40 = {5'd0, _zz_selectReadFifo_0_41};
  assign _zz_selectReadFifo_0_42 = (selectReadFifo_0 + _zz_selectReadFifo_0_43);
  assign _zz_selectReadFifo_0_43 = (3'b111 * bReg);
  assign _zz_selectReadFifo_0_45 = 1'b1;
  assign _zz_selectReadFifo_0_44 = {5'd0, _zz_selectReadFifo_0_45};
  assign _zz_when_ArraySlice_l165_208 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_208_1);
  assign _zz_when_ArraySlice_l165_208_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_208_1 = {3'd0, _zz_when_ArraySlice_l165_208_2};
  assign _zz_when_ArraySlice_l166_208 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_208_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_208_3);
  assign _zz_when_ArraySlice_l166_208_1 = {1'd0, _zz_when_ArraySlice_l166_208_2};
  assign _zz_when_ArraySlice_l166_208_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_208_4);
  assign _zz_when_ArraySlice_l166_208_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_208_4 = {3'd0, _zz_when_ArraySlice_l166_208_5};
  assign _zz__zz_when_ArraySlice_l112_208 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_208 = (_zz_when_ArraySlice_l113_208_1 - _zz_when_ArraySlice_l113_208_4);
  assign _zz_when_ArraySlice_l113_208_1 = (_zz_when_ArraySlice_l113_208_2 + _zz_when_ArraySlice_l113_208_3);
  assign _zz_when_ArraySlice_l113_208_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_208_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_208_4 = {1'd0, _zz_when_ArraySlice_l112_208};
  assign _zz__zz_when_ArraySlice_l173_208 = (_zz__zz_when_ArraySlice_l173_208_1 + _zz__zz_when_ArraySlice_l173_208_2);
  assign _zz__zz_when_ArraySlice_l173_208_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_208_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_208_3 = {1'd0, _zz_when_ArraySlice_l112_208};
  assign _zz_when_ArraySlice_l118_208_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_208 = _zz_when_ArraySlice_l118_208_1[5:0];
  assign _zz_when_ArraySlice_l173_208_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_208_2 = (_zz_when_ArraySlice_l173_208_3 + _zz_when_ArraySlice_l173_208_8);
  assign _zz_when_ArraySlice_l173_208_3 = (_zz_when_ArraySlice_l173_208 - _zz_when_ArraySlice_l173_208_4);
  assign _zz_when_ArraySlice_l173_208_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_208_6);
  assign _zz_when_ArraySlice_l173_208_4 = {1'd0, _zz_when_ArraySlice_l173_208_5};
  assign _zz_when_ArraySlice_l173_208_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_208_6 = {3'd0, _zz_when_ArraySlice_l173_208_7};
  assign _zz_when_ArraySlice_l173_208_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_209 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_209_1);
  assign _zz_when_ArraySlice_l165_209_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_209_1 = {2'd0, _zz_when_ArraySlice_l165_209_2};
  assign _zz_when_ArraySlice_l166_209 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_209_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_209_2);
  assign _zz_when_ArraySlice_l166_209_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_209_3);
  assign _zz_when_ArraySlice_l166_209_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_209_3 = {2'd0, _zz_when_ArraySlice_l166_209_4};
  assign _zz__zz_when_ArraySlice_l112_209 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_209 = (_zz_when_ArraySlice_l113_209_1 - _zz_when_ArraySlice_l113_209_4);
  assign _zz_when_ArraySlice_l113_209_1 = (_zz_when_ArraySlice_l113_209_2 + _zz_when_ArraySlice_l113_209_3);
  assign _zz_when_ArraySlice_l113_209_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_209_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_209_4 = {1'd0, _zz_when_ArraySlice_l112_209};
  assign _zz__zz_when_ArraySlice_l173_209 = (_zz__zz_when_ArraySlice_l173_209_1 + _zz__zz_when_ArraySlice_l173_209_2);
  assign _zz__zz_when_ArraySlice_l173_209_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_209_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_209_3 = {1'd0, _zz_when_ArraySlice_l112_209};
  assign _zz_when_ArraySlice_l118_209_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_209 = _zz_when_ArraySlice_l118_209_1[5:0];
  assign _zz_when_ArraySlice_l173_209_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_209_1 = {1'd0, _zz_when_ArraySlice_l173_209_2};
  assign _zz_when_ArraySlice_l173_209_3 = (_zz_when_ArraySlice_l173_209_4 + _zz_when_ArraySlice_l173_209_9);
  assign _zz_when_ArraySlice_l173_209_4 = (_zz_when_ArraySlice_l173_209 - _zz_when_ArraySlice_l173_209_5);
  assign _zz_when_ArraySlice_l173_209_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_209_7);
  assign _zz_when_ArraySlice_l173_209_5 = {1'd0, _zz_when_ArraySlice_l173_209_6};
  assign _zz_when_ArraySlice_l173_209_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_209_7 = {2'd0, _zz_when_ArraySlice_l173_209_8};
  assign _zz_when_ArraySlice_l173_209_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_210 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_210_1);
  assign _zz_when_ArraySlice_l165_210_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_210_1 = {1'd0, _zz_when_ArraySlice_l165_210_2};
  assign _zz_when_ArraySlice_l166_210 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_210_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_210_2);
  assign _zz_when_ArraySlice_l166_210_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_210_3);
  assign _zz_when_ArraySlice_l166_210_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_210_3 = {1'd0, _zz_when_ArraySlice_l166_210_4};
  assign _zz__zz_when_ArraySlice_l112_210 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_210 = (_zz_when_ArraySlice_l113_210_1 - _zz_when_ArraySlice_l113_210_4);
  assign _zz_when_ArraySlice_l113_210_1 = (_zz_when_ArraySlice_l113_210_2 + _zz_when_ArraySlice_l113_210_3);
  assign _zz_when_ArraySlice_l113_210_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_210_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_210_4 = {1'd0, _zz_when_ArraySlice_l112_210};
  assign _zz__zz_when_ArraySlice_l173_210 = (_zz__zz_when_ArraySlice_l173_210_1 + _zz__zz_when_ArraySlice_l173_210_2);
  assign _zz__zz_when_ArraySlice_l173_210_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_210_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_210_3 = {1'd0, _zz_when_ArraySlice_l112_210};
  assign _zz_when_ArraySlice_l118_210_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_210 = _zz_when_ArraySlice_l118_210_1[5:0];
  assign _zz_when_ArraySlice_l173_210_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_210_1 = {1'd0, _zz_when_ArraySlice_l173_210_2};
  assign _zz_when_ArraySlice_l173_210_3 = (_zz_when_ArraySlice_l173_210_4 + _zz_when_ArraySlice_l173_210_9);
  assign _zz_when_ArraySlice_l173_210_4 = (_zz_when_ArraySlice_l173_210 - _zz_when_ArraySlice_l173_210_5);
  assign _zz_when_ArraySlice_l173_210_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_210_7);
  assign _zz_when_ArraySlice_l173_210_5 = {1'd0, _zz_when_ArraySlice_l173_210_6};
  assign _zz_when_ArraySlice_l173_210_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_210_7 = {1'd0, _zz_when_ArraySlice_l173_210_8};
  assign _zz_when_ArraySlice_l173_210_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_211 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_211_1);
  assign _zz_when_ArraySlice_l165_211_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_211_1 = {1'd0, _zz_when_ArraySlice_l165_211_2};
  assign _zz_when_ArraySlice_l166_211 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_211_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_211_2);
  assign _zz_when_ArraySlice_l166_211_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_211_3);
  assign _zz_when_ArraySlice_l166_211_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_211_3 = {1'd0, _zz_when_ArraySlice_l166_211_4};
  assign _zz__zz_when_ArraySlice_l112_211 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_211 = (_zz_when_ArraySlice_l113_211_1 - _zz_when_ArraySlice_l113_211_4);
  assign _zz_when_ArraySlice_l113_211_1 = (_zz_when_ArraySlice_l113_211_2 + _zz_when_ArraySlice_l113_211_3);
  assign _zz_when_ArraySlice_l113_211_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_211_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_211_4 = {1'd0, _zz_when_ArraySlice_l112_211};
  assign _zz__zz_when_ArraySlice_l173_211 = (_zz__zz_when_ArraySlice_l173_211_1 + _zz__zz_when_ArraySlice_l173_211_2);
  assign _zz__zz_when_ArraySlice_l173_211_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_211_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_211_3 = {1'd0, _zz_when_ArraySlice_l112_211};
  assign _zz_when_ArraySlice_l118_211_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_211 = _zz_when_ArraySlice_l118_211_1[5:0];
  assign _zz_when_ArraySlice_l173_211_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_211_1 = {1'd0, _zz_when_ArraySlice_l173_211_2};
  assign _zz_when_ArraySlice_l173_211_3 = (_zz_when_ArraySlice_l173_211_4 + _zz_when_ArraySlice_l173_211_9);
  assign _zz_when_ArraySlice_l173_211_4 = (_zz_when_ArraySlice_l173_211 - _zz_when_ArraySlice_l173_211_5);
  assign _zz_when_ArraySlice_l173_211_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_211_7);
  assign _zz_when_ArraySlice_l173_211_5 = {1'd0, _zz_when_ArraySlice_l173_211_6};
  assign _zz_when_ArraySlice_l173_211_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_211_7 = {1'd0, _zz_when_ArraySlice_l173_211_8};
  assign _zz_when_ArraySlice_l173_211_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_212 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_212_1);
  assign _zz_when_ArraySlice_l165_212_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_212 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_212_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_212_2);
  assign _zz_when_ArraySlice_l166_212_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_212_3);
  assign _zz_when_ArraySlice_l166_212_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_212 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_212 = (_zz_when_ArraySlice_l113_212_1 - _zz_when_ArraySlice_l113_212_4);
  assign _zz_when_ArraySlice_l113_212_1 = (_zz_when_ArraySlice_l113_212_2 + _zz_when_ArraySlice_l113_212_3);
  assign _zz_when_ArraySlice_l113_212_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_212_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_212_4 = {1'd0, _zz_when_ArraySlice_l112_212};
  assign _zz__zz_when_ArraySlice_l173_212 = (_zz__zz_when_ArraySlice_l173_212_1 + _zz__zz_when_ArraySlice_l173_212_2);
  assign _zz__zz_when_ArraySlice_l173_212_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_212_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_212_3 = {1'd0, _zz_when_ArraySlice_l112_212};
  assign _zz_when_ArraySlice_l118_212_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_212 = _zz_when_ArraySlice_l118_212_1[5:0];
  assign _zz_when_ArraySlice_l173_212_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_212_1 = {1'd0, _zz_when_ArraySlice_l173_212_2};
  assign _zz_when_ArraySlice_l173_212_3 = (_zz_when_ArraySlice_l173_212_4 + _zz_when_ArraySlice_l173_212_8);
  assign _zz_when_ArraySlice_l173_212_4 = (_zz_when_ArraySlice_l173_212 - _zz_when_ArraySlice_l173_212_5);
  assign _zz_when_ArraySlice_l173_212_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_212_7);
  assign _zz_when_ArraySlice_l173_212_5 = {1'd0, _zz_when_ArraySlice_l173_212_6};
  assign _zz_when_ArraySlice_l173_212_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_212_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_213 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_213_1);
  assign _zz_when_ArraySlice_l165_213_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_213_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_213 = {1'd0, _zz_when_ArraySlice_l166_213_1};
  assign _zz_when_ArraySlice_l166_213_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_213_3);
  assign _zz_when_ArraySlice_l166_213_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_213_4);
  assign _zz_when_ArraySlice_l166_213_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_213 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_213 = (_zz_when_ArraySlice_l113_213_1 - _zz_when_ArraySlice_l113_213_4);
  assign _zz_when_ArraySlice_l113_213_1 = (_zz_when_ArraySlice_l113_213_2 + _zz_when_ArraySlice_l113_213_3);
  assign _zz_when_ArraySlice_l113_213_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_213_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_213_4 = {1'd0, _zz_when_ArraySlice_l112_213};
  assign _zz__zz_when_ArraySlice_l173_213 = (_zz__zz_when_ArraySlice_l173_213_1 + _zz__zz_when_ArraySlice_l173_213_2);
  assign _zz__zz_when_ArraySlice_l173_213_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_213_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_213_3 = {1'd0, _zz_when_ArraySlice_l112_213};
  assign _zz_when_ArraySlice_l118_213_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_213 = _zz_when_ArraySlice_l118_213_1[5:0];
  assign _zz_when_ArraySlice_l173_213_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_213_1 = {2'd0, _zz_when_ArraySlice_l173_213_2};
  assign _zz_when_ArraySlice_l173_213_3 = (_zz_when_ArraySlice_l173_213_4 + _zz_when_ArraySlice_l173_213_8);
  assign _zz_when_ArraySlice_l173_213_4 = (_zz_when_ArraySlice_l173_213 - _zz_when_ArraySlice_l173_213_5);
  assign _zz_when_ArraySlice_l173_213_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_213_7);
  assign _zz_when_ArraySlice_l173_213_5 = {1'd0, _zz_when_ArraySlice_l173_213_6};
  assign _zz_when_ArraySlice_l173_213_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_213_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_214 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_214_1);
  assign _zz_when_ArraySlice_l165_214_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_214_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_214 = {1'd0, _zz_when_ArraySlice_l166_214_1};
  assign _zz_when_ArraySlice_l166_214_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_214_3);
  assign _zz_when_ArraySlice_l166_214_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_214_4);
  assign _zz_when_ArraySlice_l166_214_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_214 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_214 = (_zz_when_ArraySlice_l113_214_1 - _zz_when_ArraySlice_l113_214_4);
  assign _zz_when_ArraySlice_l113_214_1 = (_zz_when_ArraySlice_l113_214_2 + _zz_when_ArraySlice_l113_214_3);
  assign _zz_when_ArraySlice_l113_214_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_214_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_214_4 = {1'd0, _zz_when_ArraySlice_l112_214};
  assign _zz__zz_when_ArraySlice_l173_214 = (_zz__zz_when_ArraySlice_l173_214_1 + _zz__zz_when_ArraySlice_l173_214_2);
  assign _zz__zz_when_ArraySlice_l173_214_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_214_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_214_3 = {1'd0, _zz_when_ArraySlice_l112_214};
  assign _zz_when_ArraySlice_l118_214_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_214 = _zz_when_ArraySlice_l118_214_1[5:0];
  assign _zz_when_ArraySlice_l173_214_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_214_1 = {2'd0, _zz_when_ArraySlice_l173_214_2};
  assign _zz_when_ArraySlice_l173_214_3 = (_zz_when_ArraySlice_l173_214_4 + _zz_when_ArraySlice_l173_214_8);
  assign _zz_when_ArraySlice_l173_214_4 = (_zz_when_ArraySlice_l173_214 - _zz_when_ArraySlice_l173_214_5);
  assign _zz_when_ArraySlice_l173_214_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_214_7);
  assign _zz_when_ArraySlice_l173_214_5 = {1'd0, _zz_when_ArraySlice_l173_214_6};
  assign _zz_when_ArraySlice_l173_214_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_214_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_215 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_215_1);
  assign _zz_when_ArraySlice_l165_215_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_215_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_215 = {2'd0, _zz_when_ArraySlice_l166_215_1};
  assign _zz_when_ArraySlice_l166_215_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_215_3);
  assign _zz_when_ArraySlice_l166_215_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_215_4);
  assign _zz_when_ArraySlice_l166_215_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_215 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_215 = (_zz_when_ArraySlice_l113_215_1 - _zz_when_ArraySlice_l113_215_4);
  assign _zz_when_ArraySlice_l113_215_1 = (_zz_when_ArraySlice_l113_215_2 + _zz_when_ArraySlice_l113_215_3);
  assign _zz_when_ArraySlice_l113_215_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_215_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_215_4 = {1'd0, _zz_when_ArraySlice_l112_215};
  assign _zz__zz_when_ArraySlice_l173_215 = (_zz__zz_when_ArraySlice_l173_215_1 + _zz__zz_when_ArraySlice_l173_215_2);
  assign _zz__zz_when_ArraySlice_l173_215_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_215_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_215_3 = {1'd0, _zz_when_ArraySlice_l112_215};
  assign _zz_when_ArraySlice_l118_215_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_215 = _zz_when_ArraySlice_l118_215_1[5:0];
  assign _zz_when_ArraySlice_l173_215_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_215_1 = {3'd0, _zz_when_ArraySlice_l173_215_2};
  assign _zz_when_ArraySlice_l173_215_3 = (_zz_when_ArraySlice_l173_215_4 + _zz_when_ArraySlice_l173_215_8);
  assign _zz_when_ArraySlice_l173_215_4 = (_zz_when_ArraySlice_l173_215 - _zz_when_ArraySlice_l173_215_5);
  assign _zz_when_ArraySlice_l173_215_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_215_7);
  assign _zz_when_ArraySlice_l173_215_5 = {1'd0, _zz_when_ArraySlice_l173_215_6};
  assign _zz_when_ArraySlice_l173_215_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_215_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l268 = (_zz_when_ArraySlice_l268_1 + _zz_when_ArraySlice_l268_6);
  assign _zz_when_ArraySlice_l268_1 = (_zz_when_ArraySlice_l268_2 + _zz_when_ArraySlice_l268_4);
  assign _zz_when_ArraySlice_l268_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l268_3);
  assign _zz_when_ArraySlice_l268_3 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l268_5 = 1'b1;
  assign _zz_when_ArraySlice_l268_4 = {5'd0, _zz_when_ArraySlice_l268_5};
  assign _zz_when_ArraySlice_l268_7 = 3'b000;
  assign _zz_when_ArraySlice_l268_6 = {3'd0, _zz_when_ArraySlice_l268_7};
  assign _zz_selectReadFifo_0_47 = 1'b1;
  assign _zz_selectReadFifo_0_46 = {5'd0, _zz_selectReadFifo_0_47};
  assign _zz_when_ArraySlice_l272 = (_zz_when_ArraySlice_l272_1 % aReg);
  assign _zz_when_ArraySlice_l272_1 = (handshakeTimes_0_value + _zz_when_ArraySlice_l272_2);
  assign _zz_when_ArraySlice_l272_3 = 1'b1;
  assign _zz_when_ArraySlice_l272_2 = {12'd0, _zz_when_ArraySlice_l272_3};
  assign _zz_when_ArraySlice_l276_1 = (selectReadFifo_0 + _zz_when_ArraySlice_l276_2);
  assign _zz_when_ArraySlice_l276_3 = 3'b000;
  assign _zz_when_ArraySlice_l276_2 = {3'd0, _zz_when_ArraySlice_l276_3};
  assign _zz_when_ArraySlice_l277_1 = (_zz_when_ArraySlice_l277_2 - _zz_when_ArraySlice_l277_3);
  assign _zz_when_ArraySlice_l277 = {7'd0, _zz_when_ArraySlice_l277_1};
  assign _zz_when_ArraySlice_l277_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l277_4 = 1'b1;
  assign _zz_when_ArraySlice_l277_3 = {5'd0, _zz_when_ArraySlice_l277_4};
  assign _zz__zz_when_ArraySlice_l94_25 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_25 = (_zz_when_ArraySlice_l95_25_1 - _zz_when_ArraySlice_l95_25_4);
  assign _zz_when_ArraySlice_l95_25_1 = (_zz_when_ArraySlice_l95_25_2 + _zz_when_ArraySlice_l95_25_3);
  assign _zz_when_ArraySlice_l95_25_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_25_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_25_4 = {1'd0, _zz_when_ArraySlice_l94_25};
  assign _zz__zz_when_ArraySlice_l279 = (_zz__zz_when_ArraySlice_l279_1 + _zz__zz_when_ArraySlice_l279_2);
  assign _zz__zz_when_ArraySlice_l279_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l279_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l279_3 = {1'd0, _zz_when_ArraySlice_l94_25};
  assign _zz_when_ArraySlice_l99_25_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_25 = _zz_when_ArraySlice_l99_25_1[5:0];
  assign _zz_when_ArraySlice_l279_8 = (outSliceNumb_0_value + _zz_when_ArraySlice_l279_9);
  assign _zz_when_ArraySlice_l279_10 = 1'b1;
  assign _zz_when_ArraySlice_l279_9 = {6'd0, _zz_when_ArraySlice_l279_10};
  assign _zz_when_ArraySlice_l279_11 = (_zz_when_ArraySlice_l279 / aReg);
  assign _zz_selectReadFifo_0_48 = (selectReadFifo_0 - _zz_selectReadFifo_0_49);
  assign _zz_selectReadFifo_0_49 = {3'd0, bReg};
  assign _zz_selectReadFifo_0_51 = 1'b1;
  assign _zz_selectReadFifo_0_50 = {5'd0, _zz_selectReadFifo_0_51};
  assign _zz_selectReadFifo_0_52 = (selectReadFifo_0 + _zz_selectReadFifo_0_53);
  assign _zz_selectReadFifo_0_53 = (3'b111 * bReg);
  assign _zz_selectReadFifo_0_55 = 1'b1;
  assign _zz_selectReadFifo_0_54 = {5'd0, _zz_selectReadFifo_0_55};
  assign _zz_when_ArraySlice_l165_216 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_216_1);
  assign _zz_when_ArraySlice_l165_216_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_216_1 = {3'd0, _zz_when_ArraySlice_l165_216_2};
  assign _zz_when_ArraySlice_l166_216 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_216_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_216_3);
  assign _zz_when_ArraySlice_l166_216_1 = {1'd0, _zz_when_ArraySlice_l166_216_2};
  assign _zz_when_ArraySlice_l166_216_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_216_4);
  assign _zz_when_ArraySlice_l166_216_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_216_4 = {3'd0, _zz_when_ArraySlice_l166_216_5};
  assign _zz__zz_when_ArraySlice_l112_216 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_216 = (_zz_when_ArraySlice_l113_216_1 - _zz_when_ArraySlice_l113_216_4);
  assign _zz_when_ArraySlice_l113_216_1 = (_zz_when_ArraySlice_l113_216_2 + _zz_when_ArraySlice_l113_216_3);
  assign _zz_when_ArraySlice_l113_216_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_216_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_216_4 = {1'd0, _zz_when_ArraySlice_l112_216};
  assign _zz__zz_when_ArraySlice_l173_216 = (_zz__zz_when_ArraySlice_l173_216_1 + _zz__zz_when_ArraySlice_l173_216_2);
  assign _zz__zz_when_ArraySlice_l173_216_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_216_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_216_3 = {1'd0, _zz_when_ArraySlice_l112_216};
  assign _zz_when_ArraySlice_l118_216_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_216 = _zz_when_ArraySlice_l118_216_1[5:0];
  assign _zz_when_ArraySlice_l173_216_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_216_2 = (_zz_when_ArraySlice_l173_216_3 + _zz_when_ArraySlice_l173_216_8);
  assign _zz_when_ArraySlice_l173_216_3 = (_zz_when_ArraySlice_l173_216 - _zz_when_ArraySlice_l173_216_4);
  assign _zz_when_ArraySlice_l173_216_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_216_6);
  assign _zz_when_ArraySlice_l173_216_4 = {1'd0, _zz_when_ArraySlice_l173_216_5};
  assign _zz_when_ArraySlice_l173_216_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_216_6 = {3'd0, _zz_when_ArraySlice_l173_216_7};
  assign _zz_when_ArraySlice_l173_216_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_217 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_217_1);
  assign _zz_when_ArraySlice_l165_217_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_217_1 = {2'd0, _zz_when_ArraySlice_l165_217_2};
  assign _zz_when_ArraySlice_l166_217 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_217_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_217_2);
  assign _zz_when_ArraySlice_l166_217_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_217_3);
  assign _zz_when_ArraySlice_l166_217_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_217_3 = {2'd0, _zz_when_ArraySlice_l166_217_4};
  assign _zz__zz_when_ArraySlice_l112_217 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_217 = (_zz_when_ArraySlice_l113_217_1 - _zz_when_ArraySlice_l113_217_4);
  assign _zz_when_ArraySlice_l113_217_1 = (_zz_when_ArraySlice_l113_217_2 + _zz_when_ArraySlice_l113_217_3);
  assign _zz_when_ArraySlice_l113_217_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_217_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_217_4 = {1'd0, _zz_when_ArraySlice_l112_217};
  assign _zz__zz_when_ArraySlice_l173_217 = (_zz__zz_when_ArraySlice_l173_217_1 + _zz__zz_when_ArraySlice_l173_217_2);
  assign _zz__zz_when_ArraySlice_l173_217_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_217_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_217_3 = {1'd0, _zz_when_ArraySlice_l112_217};
  assign _zz_when_ArraySlice_l118_217_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_217 = _zz_when_ArraySlice_l118_217_1[5:0];
  assign _zz_when_ArraySlice_l173_217_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_217_1 = {1'd0, _zz_when_ArraySlice_l173_217_2};
  assign _zz_when_ArraySlice_l173_217_3 = (_zz_when_ArraySlice_l173_217_4 + _zz_when_ArraySlice_l173_217_9);
  assign _zz_when_ArraySlice_l173_217_4 = (_zz_when_ArraySlice_l173_217 - _zz_when_ArraySlice_l173_217_5);
  assign _zz_when_ArraySlice_l173_217_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_217_7);
  assign _zz_when_ArraySlice_l173_217_5 = {1'd0, _zz_when_ArraySlice_l173_217_6};
  assign _zz_when_ArraySlice_l173_217_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_217_7 = {2'd0, _zz_when_ArraySlice_l173_217_8};
  assign _zz_when_ArraySlice_l173_217_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_218 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_218_1);
  assign _zz_when_ArraySlice_l165_218_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_218_1 = {1'd0, _zz_when_ArraySlice_l165_218_2};
  assign _zz_when_ArraySlice_l166_218 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_218_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_218_2);
  assign _zz_when_ArraySlice_l166_218_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_218_3);
  assign _zz_when_ArraySlice_l166_218_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_218_3 = {1'd0, _zz_when_ArraySlice_l166_218_4};
  assign _zz__zz_when_ArraySlice_l112_218 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_218 = (_zz_when_ArraySlice_l113_218_1 - _zz_when_ArraySlice_l113_218_4);
  assign _zz_when_ArraySlice_l113_218_1 = (_zz_when_ArraySlice_l113_218_2 + _zz_when_ArraySlice_l113_218_3);
  assign _zz_when_ArraySlice_l113_218_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_218_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_218_4 = {1'd0, _zz_when_ArraySlice_l112_218};
  assign _zz__zz_when_ArraySlice_l173_218 = (_zz__zz_when_ArraySlice_l173_218_1 + _zz__zz_when_ArraySlice_l173_218_2);
  assign _zz__zz_when_ArraySlice_l173_218_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_218_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_218_3 = {1'd0, _zz_when_ArraySlice_l112_218};
  assign _zz_when_ArraySlice_l118_218_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_218 = _zz_when_ArraySlice_l118_218_1[5:0];
  assign _zz_when_ArraySlice_l173_218_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_218_1 = {1'd0, _zz_when_ArraySlice_l173_218_2};
  assign _zz_when_ArraySlice_l173_218_3 = (_zz_when_ArraySlice_l173_218_4 + _zz_when_ArraySlice_l173_218_9);
  assign _zz_when_ArraySlice_l173_218_4 = (_zz_when_ArraySlice_l173_218 - _zz_when_ArraySlice_l173_218_5);
  assign _zz_when_ArraySlice_l173_218_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_218_7);
  assign _zz_when_ArraySlice_l173_218_5 = {1'd0, _zz_when_ArraySlice_l173_218_6};
  assign _zz_when_ArraySlice_l173_218_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_218_7 = {1'd0, _zz_when_ArraySlice_l173_218_8};
  assign _zz_when_ArraySlice_l173_218_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_219 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_219_1);
  assign _zz_when_ArraySlice_l165_219_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_219_1 = {1'd0, _zz_when_ArraySlice_l165_219_2};
  assign _zz_when_ArraySlice_l166_219 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_219_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_219_2);
  assign _zz_when_ArraySlice_l166_219_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_219_3);
  assign _zz_when_ArraySlice_l166_219_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_219_3 = {1'd0, _zz_when_ArraySlice_l166_219_4};
  assign _zz__zz_when_ArraySlice_l112_219 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_219 = (_zz_when_ArraySlice_l113_219_1 - _zz_when_ArraySlice_l113_219_4);
  assign _zz_when_ArraySlice_l113_219_1 = (_zz_when_ArraySlice_l113_219_2 + _zz_when_ArraySlice_l113_219_3);
  assign _zz_when_ArraySlice_l113_219_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_219_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_219_4 = {1'd0, _zz_when_ArraySlice_l112_219};
  assign _zz__zz_when_ArraySlice_l173_219 = (_zz__zz_when_ArraySlice_l173_219_1 + _zz__zz_when_ArraySlice_l173_219_2);
  assign _zz__zz_when_ArraySlice_l173_219_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_219_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_219_3 = {1'd0, _zz_when_ArraySlice_l112_219};
  assign _zz_when_ArraySlice_l118_219_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_219 = _zz_when_ArraySlice_l118_219_1[5:0];
  assign _zz_when_ArraySlice_l173_219_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_219_1 = {1'd0, _zz_when_ArraySlice_l173_219_2};
  assign _zz_when_ArraySlice_l173_219_3 = (_zz_when_ArraySlice_l173_219_4 + _zz_when_ArraySlice_l173_219_9);
  assign _zz_when_ArraySlice_l173_219_4 = (_zz_when_ArraySlice_l173_219 - _zz_when_ArraySlice_l173_219_5);
  assign _zz_when_ArraySlice_l173_219_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_219_7);
  assign _zz_when_ArraySlice_l173_219_5 = {1'd0, _zz_when_ArraySlice_l173_219_6};
  assign _zz_when_ArraySlice_l173_219_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_219_7 = {1'd0, _zz_when_ArraySlice_l173_219_8};
  assign _zz_when_ArraySlice_l173_219_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_220 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_220_1);
  assign _zz_when_ArraySlice_l165_220_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_220 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_220_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_220_2);
  assign _zz_when_ArraySlice_l166_220_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_220_3);
  assign _zz_when_ArraySlice_l166_220_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_220 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_220 = (_zz_when_ArraySlice_l113_220_1 - _zz_when_ArraySlice_l113_220_4);
  assign _zz_when_ArraySlice_l113_220_1 = (_zz_when_ArraySlice_l113_220_2 + _zz_when_ArraySlice_l113_220_3);
  assign _zz_when_ArraySlice_l113_220_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_220_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_220_4 = {1'd0, _zz_when_ArraySlice_l112_220};
  assign _zz__zz_when_ArraySlice_l173_220 = (_zz__zz_when_ArraySlice_l173_220_1 + _zz__zz_when_ArraySlice_l173_220_2);
  assign _zz__zz_when_ArraySlice_l173_220_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_220_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_220_3 = {1'd0, _zz_when_ArraySlice_l112_220};
  assign _zz_when_ArraySlice_l118_220_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_220 = _zz_when_ArraySlice_l118_220_1[5:0];
  assign _zz_when_ArraySlice_l173_220_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_220_1 = {1'd0, _zz_when_ArraySlice_l173_220_2};
  assign _zz_when_ArraySlice_l173_220_3 = (_zz_when_ArraySlice_l173_220_4 + _zz_when_ArraySlice_l173_220_8);
  assign _zz_when_ArraySlice_l173_220_4 = (_zz_when_ArraySlice_l173_220 - _zz_when_ArraySlice_l173_220_5);
  assign _zz_when_ArraySlice_l173_220_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_220_7);
  assign _zz_when_ArraySlice_l173_220_5 = {1'd0, _zz_when_ArraySlice_l173_220_6};
  assign _zz_when_ArraySlice_l173_220_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_220_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_221 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_221_1);
  assign _zz_when_ArraySlice_l165_221_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_221_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_221 = {1'd0, _zz_when_ArraySlice_l166_221_1};
  assign _zz_when_ArraySlice_l166_221_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_221_3);
  assign _zz_when_ArraySlice_l166_221_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_221_4);
  assign _zz_when_ArraySlice_l166_221_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_221 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_221 = (_zz_when_ArraySlice_l113_221_1 - _zz_when_ArraySlice_l113_221_4);
  assign _zz_when_ArraySlice_l113_221_1 = (_zz_when_ArraySlice_l113_221_2 + _zz_when_ArraySlice_l113_221_3);
  assign _zz_when_ArraySlice_l113_221_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_221_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_221_4 = {1'd0, _zz_when_ArraySlice_l112_221};
  assign _zz__zz_when_ArraySlice_l173_221 = (_zz__zz_when_ArraySlice_l173_221_1 + _zz__zz_when_ArraySlice_l173_221_2);
  assign _zz__zz_when_ArraySlice_l173_221_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_221_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_221_3 = {1'd0, _zz_when_ArraySlice_l112_221};
  assign _zz_when_ArraySlice_l118_221_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_221 = _zz_when_ArraySlice_l118_221_1[5:0];
  assign _zz_when_ArraySlice_l173_221_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_221_1 = {2'd0, _zz_when_ArraySlice_l173_221_2};
  assign _zz_when_ArraySlice_l173_221_3 = (_zz_when_ArraySlice_l173_221_4 + _zz_when_ArraySlice_l173_221_8);
  assign _zz_when_ArraySlice_l173_221_4 = (_zz_when_ArraySlice_l173_221 - _zz_when_ArraySlice_l173_221_5);
  assign _zz_when_ArraySlice_l173_221_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_221_7);
  assign _zz_when_ArraySlice_l173_221_5 = {1'd0, _zz_when_ArraySlice_l173_221_6};
  assign _zz_when_ArraySlice_l173_221_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_221_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_222 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_222_1);
  assign _zz_when_ArraySlice_l165_222_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_222_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_222 = {1'd0, _zz_when_ArraySlice_l166_222_1};
  assign _zz_when_ArraySlice_l166_222_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_222_3);
  assign _zz_when_ArraySlice_l166_222_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_222_4);
  assign _zz_when_ArraySlice_l166_222_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_222 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_222 = (_zz_when_ArraySlice_l113_222_1 - _zz_when_ArraySlice_l113_222_4);
  assign _zz_when_ArraySlice_l113_222_1 = (_zz_when_ArraySlice_l113_222_2 + _zz_when_ArraySlice_l113_222_3);
  assign _zz_when_ArraySlice_l113_222_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_222_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_222_4 = {1'd0, _zz_when_ArraySlice_l112_222};
  assign _zz__zz_when_ArraySlice_l173_222 = (_zz__zz_when_ArraySlice_l173_222_1 + _zz__zz_when_ArraySlice_l173_222_2);
  assign _zz__zz_when_ArraySlice_l173_222_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_222_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_222_3 = {1'd0, _zz_when_ArraySlice_l112_222};
  assign _zz_when_ArraySlice_l118_222_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_222 = _zz_when_ArraySlice_l118_222_1[5:0];
  assign _zz_when_ArraySlice_l173_222_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_222_1 = {2'd0, _zz_when_ArraySlice_l173_222_2};
  assign _zz_when_ArraySlice_l173_222_3 = (_zz_when_ArraySlice_l173_222_4 + _zz_when_ArraySlice_l173_222_8);
  assign _zz_when_ArraySlice_l173_222_4 = (_zz_when_ArraySlice_l173_222 - _zz_when_ArraySlice_l173_222_5);
  assign _zz_when_ArraySlice_l173_222_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_222_7);
  assign _zz_when_ArraySlice_l173_222_5 = {1'd0, _zz_when_ArraySlice_l173_222_6};
  assign _zz_when_ArraySlice_l173_222_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_222_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_223 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_223_1);
  assign _zz_when_ArraySlice_l165_223_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_223_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_223 = {2'd0, _zz_when_ArraySlice_l166_223_1};
  assign _zz_when_ArraySlice_l166_223_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_223_3);
  assign _zz_when_ArraySlice_l166_223_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_223_4);
  assign _zz_when_ArraySlice_l166_223_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_223 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_223 = (_zz_when_ArraySlice_l113_223_1 - _zz_when_ArraySlice_l113_223_4);
  assign _zz_when_ArraySlice_l113_223_1 = (_zz_when_ArraySlice_l113_223_2 + _zz_when_ArraySlice_l113_223_3);
  assign _zz_when_ArraySlice_l113_223_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_223_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_223_4 = {1'd0, _zz_when_ArraySlice_l112_223};
  assign _zz__zz_when_ArraySlice_l173_223 = (_zz__zz_when_ArraySlice_l173_223_1 + _zz__zz_when_ArraySlice_l173_223_2);
  assign _zz__zz_when_ArraySlice_l173_223_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_223_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_223_3 = {1'd0, _zz_when_ArraySlice_l112_223};
  assign _zz_when_ArraySlice_l118_223_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_223 = _zz_when_ArraySlice_l118_223_1[5:0];
  assign _zz_when_ArraySlice_l173_223_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_223_1 = {3'd0, _zz_when_ArraySlice_l173_223_2};
  assign _zz_when_ArraySlice_l173_223_3 = (_zz_when_ArraySlice_l173_223_4 + _zz_when_ArraySlice_l173_223_8);
  assign _zz_when_ArraySlice_l173_223_4 = (_zz_when_ArraySlice_l173_223 - _zz_when_ArraySlice_l173_223_5);
  assign _zz_when_ArraySlice_l173_223_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_223_7);
  assign _zz_when_ArraySlice_l173_223_5 = {1'd0, _zz_when_ArraySlice_l173_223_6};
  assign _zz_when_ArraySlice_l173_223_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_223_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l288 = (_zz_when_ArraySlice_l288_1 + _zz_when_ArraySlice_l288_6);
  assign _zz_when_ArraySlice_l288_1 = (_zz_when_ArraySlice_l288_2 + _zz_when_ArraySlice_l288_4);
  assign _zz_when_ArraySlice_l288_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l288_3);
  assign _zz_when_ArraySlice_l288_3 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_5 = 1'b1;
  assign _zz_when_ArraySlice_l288_4 = {5'd0, _zz_when_ArraySlice_l288_5};
  assign _zz_when_ArraySlice_l288_7 = 3'b000;
  assign _zz_when_ArraySlice_l288_6 = {3'd0, _zz_when_ArraySlice_l288_7};
  assign _zz_selectReadFifo_0_57 = 1'b1;
  assign _zz_selectReadFifo_0_56 = {5'd0, _zz_selectReadFifo_0_57};
  assign _zz_when_ArraySlice_l292 = (_zz_when_ArraySlice_l292_1 % aReg);
  assign _zz_when_ArraySlice_l292_1 = (handshakeTimes_0_value + _zz_when_ArraySlice_l292_2);
  assign _zz_when_ArraySlice_l292_3 = 1'b1;
  assign _zz_when_ArraySlice_l292_2 = {12'd0, _zz_when_ArraySlice_l292_3};
  assign _zz_when_ArraySlice_l303_1 = (_zz_when_ArraySlice_l303_2 - _zz_when_ArraySlice_l303_3);
  assign _zz_when_ArraySlice_l303 = {7'd0, _zz_when_ArraySlice_l303_1};
  assign _zz_when_ArraySlice_l303_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l303_4 = 1'b1;
  assign _zz_when_ArraySlice_l303_3 = {5'd0, _zz_when_ArraySlice_l303_4};
  assign _zz__zz_when_ArraySlice_l94_26 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_26 = (_zz_when_ArraySlice_l95_26_1 - _zz_when_ArraySlice_l95_26_4);
  assign _zz_when_ArraySlice_l95_26_1 = (_zz_when_ArraySlice_l95_26_2 + _zz_when_ArraySlice_l95_26_3);
  assign _zz_when_ArraySlice_l95_26_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_26_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_26_4 = {1'd0, _zz_when_ArraySlice_l94_26};
  assign _zz__zz_when_ArraySlice_l304 = (_zz__zz_when_ArraySlice_l304_1 + _zz__zz_when_ArraySlice_l304_2);
  assign _zz__zz_when_ArraySlice_l304_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l304_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l304_3 = {1'd0, _zz_when_ArraySlice_l94_26};
  assign _zz_when_ArraySlice_l99_26_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_26 = _zz_when_ArraySlice_l99_26_1[5:0];
  assign _zz_when_ArraySlice_l304_8 = (outSliceNumb_0_value + _zz_when_ArraySlice_l304_9);
  assign _zz_when_ArraySlice_l304_10 = 1'b1;
  assign _zz_when_ArraySlice_l304_9 = {6'd0, _zz_when_ArraySlice_l304_10};
  assign _zz_when_ArraySlice_l304_11 = (_zz_when_ArraySlice_l304 / aReg);
  assign _zz_selectReadFifo_0_58 = (selectReadFifo_0 - _zz_selectReadFifo_0_59);
  assign _zz_selectReadFifo_0_59 = {3'd0, bReg};
  assign _zz_selectReadFifo_0_61 = 1'b1;
  assign _zz_selectReadFifo_0_60 = {5'd0, _zz_selectReadFifo_0_61};
  assign _zz_when_ArraySlice_l165_224 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_224_1);
  assign _zz_when_ArraySlice_l165_224_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_224_1 = {3'd0, _zz_when_ArraySlice_l165_224_2};
  assign _zz_when_ArraySlice_l166_224 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_224_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_224_3);
  assign _zz_when_ArraySlice_l166_224_1 = {1'd0, _zz_when_ArraySlice_l166_224_2};
  assign _zz_when_ArraySlice_l166_224_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_224_4);
  assign _zz_when_ArraySlice_l166_224_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_224_4 = {3'd0, _zz_when_ArraySlice_l166_224_5};
  assign _zz__zz_when_ArraySlice_l112_224 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_224 = (_zz_when_ArraySlice_l113_224_1 - _zz_when_ArraySlice_l113_224_4);
  assign _zz_when_ArraySlice_l113_224_1 = (_zz_when_ArraySlice_l113_224_2 + _zz_when_ArraySlice_l113_224_3);
  assign _zz_when_ArraySlice_l113_224_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_224_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_224_4 = {1'd0, _zz_when_ArraySlice_l112_224};
  assign _zz__zz_when_ArraySlice_l173_224 = (_zz__zz_when_ArraySlice_l173_224_1 + _zz__zz_when_ArraySlice_l173_224_2);
  assign _zz__zz_when_ArraySlice_l173_224_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_224_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_224_3 = {1'd0, _zz_when_ArraySlice_l112_224};
  assign _zz_when_ArraySlice_l118_224_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_224 = _zz_when_ArraySlice_l118_224_1[5:0];
  assign _zz_when_ArraySlice_l173_224_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_224_2 = (_zz_when_ArraySlice_l173_224_3 + _zz_when_ArraySlice_l173_224_8);
  assign _zz_when_ArraySlice_l173_224_3 = (_zz_when_ArraySlice_l173_224 - _zz_when_ArraySlice_l173_224_4);
  assign _zz_when_ArraySlice_l173_224_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_224_6);
  assign _zz_when_ArraySlice_l173_224_4 = {1'd0, _zz_when_ArraySlice_l173_224_5};
  assign _zz_when_ArraySlice_l173_224_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_224_6 = {3'd0, _zz_when_ArraySlice_l173_224_7};
  assign _zz_when_ArraySlice_l173_224_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_225 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_225_1);
  assign _zz_when_ArraySlice_l165_225_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_225_1 = {2'd0, _zz_when_ArraySlice_l165_225_2};
  assign _zz_when_ArraySlice_l166_225 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_225_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_225_2);
  assign _zz_when_ArraySlice_l166_225_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_225_3);
  assign _zz_when_ArraySlice_l166_225_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_225_3 = {2'd0, _zz_when_ArraySlice_l166_225_4};
  assign _zz__zz_when_ArraySlice_l112_225 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_225 = (_zz_when_ArraySlice_l113_225_1 - _zz_when_ArraySlice_l113_225_4);
  assign _zz_when_ArraySlice_l113_225_1 = (_zz_when_ArraySlice_l113_225_2 + _zz_when_ArraySlice_l113_225_3);
  assign _zz_when_ArraySlice_l113_225_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_225_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_225_4 = {1'd0, _zz_when_ArraySlice_l112_225};
  assign _zz__zz_when_ArraySlice_l173_225 = (_zz__zz_when_ArraySlice_l173_225_1 + _zz__zz_when_ArraySlice_l173_225_2);
  assign _zz__zz_when_ArraySlice_l173_225_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_225_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_225_3 = {1'd0, _zz_when_ArraySlice_l112_225};
  assign _zz_when_ArraySlice_l118_225_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_225 = _zz_when_ArraySlice_l118_225_1[5:0];
  assign _zz_when_ArraySlice_l173_225_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_225_1 = {1'd0, _zz_when_ArraySlice_l173_225_2};
  assign _zz_when_ArraySlice_l173_225_3 = (_zz_when_ArraySlice_l173_225_4 + _zz_when_ArraySlice_l173_225_9);
  assign _zz_when_ArraySlice_l173_225_4 = (_zz_when_ArraySlice_l173_225 - _zz_when_ArraySlice_l173_225_5);
  assign _zz_when_ArraySlice_l173_225_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_225_7);
  assign _zz_when_ArraySlice_l173_225_5 = {1'd0, _zz_when_ArraySlice_l173_225_6};
  assign _zz_when_ArraySlice_l173_225_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_225_7 = {2'd0, _zz_when_ArraySlice_l173_225_8};
  assign _zz_when_ArraySlice_l173_225_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_226 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_226_1);
  assign _zz_when_ArraySlice_l165_226_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_226_1 = {1'd0, _zz_when_ArraySlice_l165_226_2};
  assign _zz_when_ArraySlice_l166_226 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_226_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_226_2);
  assign _zz_when_ArraySlice_l166_226_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_226_3);
  assign _zz_when_ArraySlice_l166_226_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_226_3 = {1'd0, _zz_when_ArraySlice_l166_226_4};
  assign _zz__zz_when_ArraySlice_l112_226 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_226 = (_zz_when_ArraySlice_l113_226_1 - _zz_when_ArraySlice_l113_226_4);
  assign _zz_when_ArraySlice_l113_226_1 = (_zz_when_ArraySlice_l113_226_2 + _zz_when_ArraySlice_l113_226_3);
  assign _zz_when_ArraySlice_l113_226_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_226_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_226_4 = {1'd0, _zz_when_ArraySlice_l112_226};
  assign _zz__zz_when_ArraySlice_l173_226 = (_zz__zz_when_ArraySlice_l173_226_1 + _zz__zz_when_ArraySlice_l173_226_2);
  assign _zz__zz_when_ArraySlice_l173_226_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_226_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_226_3 = {1'd0, _zz_when_ArraySlice_l112_226};
  assign _zz_when_ArraySlice_l118_226_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_226 = _zz_when_ArraySlice_l118_226_1[5:0];
  assign _zz_when_ArraySlice_l173_226_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_226_1 = {1'd0, _zz_when_ArraySlice_l173_226_2};
  assign _zz_when_ArraySlice_l173_226_3 = (_zz_when_ArraySlice_l173_226_4 + _zz_when_ArraySlice_l173_226_9);
  assign _zz_when_ArraySlice_l173_226_4 = (_zz_when_ArraySlice_l173_226 - _zz_when_ArraySlice_l173_226_5);
  assign _zz_when_ArraySlice_l173_226_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_226_7);
  assign _zz_when_ArraySlice_l173_226_5 = {1'd0, _zz_when_ArraySlice_l173_226_6};
  assign _zz_when_ArraySlice_l173_226_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_226_7 = {1'd0, _zz_when_ArraySlice_l173_226_8};
  assign _zz_when_ArraySlice_l173_226_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_227 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_227_1);
  assign _zz_when_ArraySlice_l165_227_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_227_1 = {1'd0, _zz_when_ArraySlice_l165_227_2};
  assign _zz_when_ArraySlice_l166_227 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_227_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_227_2);
  assign _zz_when_ArraySlice_l166_227_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_227_3);
  assign _zz_when_ArraySlice_l166_227_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_227_3 = {1'd0, _zz_when_ArraySlice_l166_227_4};
  assign _zz__zz_when_ArraySlice_l112_227 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_227 = (_zz_when_ArraySlice_l113_227_1 - _zz_when_ArraySlice_l113_227_4);
  assign _zz_when_ArraySlice_l113_227_1 = (_zz_when_ArraySlice_l113_227_2 + _zz_when_ArraySlice_l113_227_3);
  assign _zz_when_ArraySlice_l113_227_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_227_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_227_4 = {1'd0, _zz_when_ArraySlice_l112_227};
  assign _zz__zz_when_ArraySlice_l173_227 = (_zz__zz_when_ArraySlice_l173_227_1 + _zz__zz_when_ArraySlice_l173_227_2);
  assign _zz__zz_when_ArraySlice_l173_227_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_227_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_227_3 = {1'd0, _zz_when_ArraySlice_l112_227};
  assign _zz_when_ArraySlice_l118_227_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_227 = _zz_when_ArraySlice_l118_227_1[5:0];
  assign _zz_when_ArraySlice_l173_227_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_227_1 = {1'd0, _zz_when_ArraySlice_l173_227_2};
  assign _zz_when_ArraySlice_l173_227_3 = (_zz_when_ArraySlice_l173_227_4 + _zz_when_ArraySlice_l173_227_9);
  assign _zz_when_ArraySlice_l173_227_4 = (_zz_when_ArraySlice_l173_227 - _zz_when_ArraySlice_l173_227_5);
  assign _zz_when_ArraySlice_l173_227_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_227_7);
  assign _zz_when_ArraySlice_l173_227_5 = {1'd0, _zz_when_ArraySlice_l173_227_6};
  assign _zz_when_ArraySlice_l173_227_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_227_7 = {1'd0, _zz_when_ArraySlice_l173_227_8};
  assign _zz_when_ArraySlice_l173_227_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_228 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_228_1);
  assign _zz_when_ArraySlice_l165_228_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_228 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_228_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_228_2);
  assign _zz_when_ArraySlice_l166_228_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_228_3);
  assign _zz_when_ArraySlice_l166_228_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_228 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_228 = (_zz_when_ArraySlice_l113_228_1 - _zz_when_ArraySlice_l113_228_4);
  assign _zz_when_ArraySlice_l113_228_1 = (_zz_when_ArraySlice_l113_228_2 + _zz_when_ArraySlice_l113_228_3);
  assign _zz_when_ArraySlice_l113_228_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_228_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_228_4 = {1'd0, _zz_when_ArraySlice_l112_228};
  assign _zz__zz_when_ArraySlice_l173_228 = (_zz__zz_when_ArraySlice_l173_228_1 + _zz__zz_when_ArraySlice_l173_228_2);
  assign _zz__zz_when_ArraySlice_l173_228_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_228_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_228_3 = {1'd0, _zz_when_ArraySlice_l112_228};
  assign _zz_when_ArraySlice_l118_228_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_228 = _zz_when_ArraySlice_l118_228_1[5:0];
  assign _zz_when_ArraySlice_l173_228_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_228_1 = {1'd0, _zz_when_ArraySlice_l173_228_2};
  assign _zz_when_ArraySlice_l173_228_3 = (_zz_when_ArraySlice_l173_228_4 + _zz_when_ArraySlice_l173_228_8);
  assign _zz_when_ArraySlice_l173_228_4 = (_zz_when_ArraySlice_l173_228 - _zz_when_ArraySlice_l173_228_5);
  assign _zz_when_ArraySlice_l173_228_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_228_7);
  assign _zz_when_ArraySlice_l173_228_5 = {1'd0, _zz_when_ArraySlice_l173_228_6};
  assign _zz_when_ArraySlice_l173_228_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_228_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_229 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_229_1);
  assign _zz_when_ArraySlice_l165_229_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_229_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_229 = {1'd0, _zz_when_ArraySlice_l166_229_1};
  assign _zz_when_ArraySlice_l166_229_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_229_3);
  assign _zz_when_ArraySlice_l166_229_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_229_4);
  assign _zz_when_ArraySlice_l166_229_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_229 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_229 = (_zz_when_ArraySlice_l113_229_1 - _zz_when_ArraySlice_l113_229_4);
  assign _zz_when_ArraySlice_l113_229_1 = (_zz_when_ArraySlice_l113_229_2 + _zz_when_ArraySlice_l113_229_3);
  assign _zz_when_ArraySlice_l113_229_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_229_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_229_4 = {1'd0, _zz_when_ArraySlice_l112_229};
  assign _zz__zz_when_ArraySlice_l173_229 = (_zz__zz_when_ArraySlice_l173_229_1 + _zz__zz_when_ArraySlice_l173_229_2);
  assign _zz__zz_when_ArraySlice_l173_229_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_229_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_229_3 = {1'd0, _zz_when_ArraySlice_l112_229};
  assign _zz_when_ArraySlice_l118_229_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_229 = _zz_when_ArraySlice_l118_229_1[5:0];
  assign _zz_when_ArraySlice_l173_229_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_229_1 = {2'd0, _zz_when_ArraySlice_l173_229_2};
  assign _zz_when_ArraySlice_l173_229_3 = (_zz_when_ArraySlice_l173_229_4 + _zz_when_ArraySlice_l173_229_8);
  assign _zz_when_ArraySlice_l173_229_4 = (_zz_when_ArraySlice_l173_229 - _zz_when_ArraySlice_l173_229_5);
  assign _zz_when_ArraySlice_l173_229_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_229_7);
  assign _zz_when_ArraySlice_l173_229_5 = {1'd0, _zz_when_ArraySlice_l173_229_6};
  assign _zz_when_ArraySlice_l173_229_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_229_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_230 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_230_1);
  assign _zz_when_ArraySlice_l165_230_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_230_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_230 = {1'd0, _zz_when_ArraySlice_l166_230_1};
  assign _zz_when_ArraySlice_l166_230_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_230_3);
  assign _zz_when_ArraySlice_l166_230_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_230_4);
  assign _zz_when_ArraySlice_l166_230_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_230 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_230 = (_zz_when_ArraySlice_l113_230_1 - _zz_when_ArraySlice_l113_230_4);
  assign _zz_when_ArraySlice_l113_230_1 = (_zz_when_ArraySlice_l113_230_2 + _zz_when_ArraySlice_l113_230_3);
  assign _zz_when_ArraySlice_l113_230_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_230_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_230_4 = {1'd0, _zz_when_ArraySlice_l112_230};
  assign _zz__zz_when_ArraySlice_l173_230 = (_zz__zz_when_ArraySlice_l173_230_1 + _zz__zz_when_ArraySlice_l173_230_2);
  assign _zz__zz_when_ArraySlice_l173_230_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_230_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_230_3 = {1'd0, _zz_when_ArraySlice_l112_230};
  assign _zz_when_ArraySlice_l118_230_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_230 = _zz_when_ArraySlice_l118_230_1[5:0];
  assign _zz_when_ArraySlice_l173_230_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_230_1 = {2'd0, _zz_when_ArraySlice_l173_230_2};
  assign _zz_when_ArraySlice_l173_230_3 = (_zz_when_ArraySlice_l173_230_4 + _zz_when_ArraySlice_l173_230_8);
  assign _zz_when_ArraySlice_l173_230_4 = (_zz_when_ArraySlice_l173_230 - _zz_when_ArraySlice_l173_230_5);
  assign _zz_when_ArraySlice_l173_230_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_230_7);
  assign _zz_when_ArraySlice_l173_230_5 = {1'd0, _zz_when_ArraySlice_l173_230_6};
  assign _zz_when_ArraySlice_l173_230_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_230_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_231 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_231_1);
  assign _zz_when_ArraySlice_l165_231_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_231_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_231 = {2'd0, _zz_when_ArraySlice_l166_231_1};
  assign _zz_when_ArraySlice_l166_231_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_231_3);
  assign _zz_when_ArraySlice_l166_231_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_231_4);
  assign _zz_when_ArraySlice_l166_231_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_231 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_231 = (_zz_when_ArraySlice_l113_231_1 - _zz_when_ArraySlice_l113_231_4);
  assign _zz_when_ArraySlice_l113_231_1 = (_zz_when_ArraySlice_l113_231_2 + _zz_when_ArraySlice_l113_231_3);
  assign _zz_when_ArraySlice_l113_231_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_231_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_231_4 = {1'd0, _zz_when_ArraySlice_l112_231};
  assign _zz__zz_when_ArraySlice_l173_231 = (_zz__zz_when_ArraySlice_l173_231_1 + _zz__zz_when_ArraySlice_l173_231_2);
  assign _zz__zz_when_ArraySlice_l173_231_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_231_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_231_3 = {1'd0, _zz_when_ArraySlice_l112_231};
  assign _zz_when_ArraySlice_l118_231_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_231 = _zz_when_ArraySlice_l118_231_1[5:0];
  assign _zz_when_ArraySlice_l173_231_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_231_1 = {3'd0, _zz_when_ArraySlice_l173_231_2};
  assign _zz_when_ArraySlice_l173_231_3 = (_zz_when_ArraySlice_l173_231_4 + _zz_when_ArraySlice_l173_231_8);
  assign _zz_when_ArraySlice_l173_231_4 = (_zz_when_ArraySlice_l173_231 - _zz_when_ArraySlice_l173_231_5);
  assign _zz_when_ArraySlice_l173_231_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_231_7);
  assign _zz_when_ArraySlice_l173_231_5 = {1'd0, _zz_when_ArraySlice_l173_231_6};
  assign _zz_when_ArraySlice_l173_231_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_231_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_0_63 = 1'b1;
  assign _zz_selectReadFifo_0_62 = {5'd0, _zz_selectReadFifo_0_63};
  assign _zz_when_ArraySlice_l315 = (_zz_when_ArraySlice_l315_1 % aReg);
  assign _zz_when_ArraySlice_l315_1 = (handshakeTimes_0_value + _zz_when_ArraySlice_l315_2);
  assign _zz_when_ArraySlice_l315_3 = 1'b1;
  assign _zz_when_ArraySlice_l315_2 = {12'd0, _zz_when_ArraySlice_l315_3};
  assign _zz_when_ArraySlice_l301 = (selectReadFifo_0 + _zz_when_ArraySlice_l301_1);
  assign _zz_when_ArraySlice_l301_2 = 3'b000;
  assign _zz_when_ArraySlice_l301_1 = {3'd0, _zz_when_ArraySlice_l301_2};
  assign _zz_when_ArraySlice_l322_1 = (_zz_when_ArraySlice_l322_2 - _zz_when_ArraySlice_l322_3);
  assign _zz_when_ArraySlice_l322 = {7'd0, _zz_when_ArraySlice_l322_1};
  assign _zz_when_ArraySlice_l322_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l322_4 = 1'b1;
  assign _zz_when_ArraySlice_l322_3 = {5'd0, _zz_when_ArraySlice_l322_4};
  assign _zz_when_ArraySlice_l240_1_1 = (selectReadFifo_1 + _zz_when_ArraySlice_l240_1_2);
  assign _zz_when_ArraySlice_l240_1_3 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l240_1_2 = {2'd0, _zz_when_ArraySlice_l240_1_3};
  assign _zz_when_ArraySlice_l241_1_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l241_1_3);
  assign _zz_when_ArraySlice_l241_1_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l241_1_3 = {2'd0, _zz_when_ArraySlice_l241_1_4};
  assign _zz__zz_outputStreamArrayData_1_valid_1_2 = (bReg * 1'b1);
  assign _zz__zz_outputStreamArrayData_1_valid_1_1 = {2'd0, _zz__zz_outputStreamArrayData_1_valid_1_2};
  assign _zz_when_ArraySlice_l247_1_2 = 1'b1;
  assign _zz_when_ArraySlice_l247_1_1 = {6'd0, _zz_when_ArraySlice_l247_1_2};
  assign _zz_when_ArraySlice_l247_1_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l247_1_5);
  assign _zz_when_ArraySlice_l247_1_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l247_1_5 = {2'd0, _zz_when_ArraySlice_l247_1_6};
  assign _zz_when_ArraySlice_l248_1_2 = (_zz_when_ArraySlice_l248_1_3 - _zz_when_ArraySlice_l248_1_4);
  assign _zz_when_ArraySlice_l248_1_1 = {7'd0, _zz_when_ArraySlice_l248_1_2};
  assign _zz_when_ArraySlice_l248_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l248_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l248_1_4 = {5'd0, _zz_when_ArraySlice_l248_1_5};
  assign _zz_selectReadFifo_1_32 = (selectReadFifo_1 - _zz_selectReadFifo_1_33);
  assign _zz_selectReadFifo_1_33 = {3'd0, bReg};
  assign _zz_selectReadFifo_1_35 = 1'b1;
  assign _zz_selectReadFifo_1_34 = {5'd0, _zz_selectReadFifo_1_35};
  assign _zz_selectReadFifo_1_37 = 1'b1;
  assign _zz_selectReadFifo_1_36 = {5'd0, _zz_selectReadFifo_1_37};
  assign _zz_when_ArraySlice_l251_1_1 = (_zz_when_ArraySlice_l251_1_2 % aReg);
  assign _zz_when_ArraySlice_l251_1_2 = (handshakeTimes_1_value + _zz_when_ArraySlice_l251_1_3);
  assign _zz_when_ArraySlice_l251_1_4 = 1'b1;
  assign _zz_when_ArraySlice_l251_1_3 = {12'd0, _zz_when_ArraySlice_l251_1_4};
  assign _zz_when_ArraySlice_l256_1_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l256_1_3);
  assign _zz_when_ArraySlice_l256_1_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l256_1_3 = {2'd0, _zz_when_ArraySlice_l256_1_4};
  assign _zz_when_ArraySlice_l256_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l256_1_5 = {6'd0, _zz_when_ArraySlice_l256_1_6};
  assign _zz_when_ArraySlice_l257_1_2 = (_zz_when_ArraySlice_l257_1_3 - _zz_when_ArraySlice_l257_1_4);
  assign _zz_when_ArraySlice_l257_1_1 = {7'd0, _zz_when_ArraySlice_l257_1_2};
  assign _zz_when_ArraySlice_l257_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l257_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l257_1_4 = {5'd0, _zz_when_ArraySlice_l257_1_5};
  assign _zz__zz_when_ArraySlice_l94_27 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_27 = (_zz_when_ArraySlice_l95_27_1 - _zz_when_ArraySlice_l95_27_4);
  assign _zz_when_ArraySlice_l95_27_1 = (_zz_when_ArraySlice_l95_27_2 + _zz_when_ArraySlice_l95_27_3);
  assign _zz_when_ArraySlice_l95_27_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_27_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_27_4 = {1'd0, _zz_when_ArraySlice_l94_27};
  assign _zz__zz_when_ArraySlice_l259_1_1 = (_zz__zz_when_ArraySlice_l259_1_2 + _zz__zz_when_ArraySlice_l259_1_3);
  assign _zz__zz_when_ArraySlice_l259_1_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l259_1_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l259_1_4 = {1'd0, _zz_when_ArraySlice_l94_27};
  assign _zz_when_ArraySlice_l99_27_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_27 = _zz_when_ArraySlice_l99_27_1[5:0];
  assign _zz_when_ArraySlice_l259_1_1 = (outSliceNumb_1_value + _zz_when_ArraySlice_l259_1_2);
  assign _zz_when_ArraySlice_l259_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l259_1_2 = {6'd0, _zz_when_ArraySlice_l259_1_3};
  assign _zz_when_ArraySlice_l259_1_4 = (_zz_when_ArraySlice_l259_1 / aReg);
  assign _zz_selectReadFifo_1_38 = (selectReadFifo_1 - _zz_selectReadFifo_1_39);
  assign _zz_selectReadFifo_1_39 = {3'd0, bReg};
  assign _zz_selectReadFifo_1_41 = 1'b1;
  assign _zz_selectReadFifo_1_40 = {5'd0, _zz_selectReadFifo_1_41};
  assign _zz_selectReadFifo_1_42 = (selectReadFifo_1 + _zz_selectReadFifo_1_43);
  assign _zz_selectReadFifo_1_43 = (3'b111 * bReg);
  assign _zz_selectReadFifo_1_45 = 1'b1;
  assign _zz_selectReadFifo_1_44 = {5'd0, _zz_selectReadFifo_1_45};
  assign _zz_when_ArraySlice_l165_232 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_232_1);
  assign _zz_when_ArraySlice_l165_232_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_232_1 = {3'd0, _zz_when_ArraySlice_l165_232_2};
  assign _zz_when_ArraySlice_l166_232 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_232_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_232_3);
  assign _zz_when_ArraySlice_l166_232_1 = {1'd0, _zz_when_ArraySlice_l166_232_2};
  assign _zz_when_ArraySlice_l166_232_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_232_4);
  assign _zz_when_ArraySlice_l166_232_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_232_4 = {3'd0, _zz_when_ArraySlice_l166_232_5};
  assign _zz__zz_when_ArraySlice_l112_232 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_232 = (_zz_when_ArraySlice_l113_232_1 - _zz_when_ArraySlice_l113_232_4);
  assign _zz_when_ArraySlice_l113_232_1 = (_zz_when_ArraySlice_l113_232_2 + _zz_when_ArraySlice_l113_232_3);
  assign _zz_when_ArraySlice_l113_232_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_232_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_232_4 = {1'd0, _zz_when_ArraySlice_l112_232};
  assign _zz__zz_when_ArraySlice_l173_232 = (_zz__zz_when_ArraySlice_l173_232_1 + _zz__zz_when_ArraySlice_l173_232_2);
  assign _zz__zz_when_ArraySlice_l173_232_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_232_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_232_3 = {1'd0, _zz_when_ArraySlice_l112_232};
  assign _zz_when_ArraySlice_l118_232_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_232 = _zz_when_ArraySlice_l118_232_1[5:0];
  assign _zz_when_ArraySlice_l173_232_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_232_2 = (_zz_when_ArraySlice_l173_232_3 + _zz_when_ArraySlice_l173_232_8);
  assign _zz_when_ArraySlice_l173_232_3 = (_zz_when_ArraySlice_l173_232 - _zz_when_ArraySlice_l173_232_4);
  assign _zz_when_ArraySlice_l173_232_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_232_6);
  assign _zz_when_ArraySlice_l173_232_4 = {1'd0, _zz_when_ArraySlice_l173_232_5};
  assign _zz_when_ArraySlice_l173_232_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_232_6 = {3'd0, _zz_when_ArraySlice_l173_232_7};
  assign _zz_when_ArraySlice_l173_232_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_233 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_233_1);
  assign _zz_when_ArraySlice_l165_233_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_233_1 = {2'd0, _zz_when_ArraySlice_l165_233_2};
  assign _zz_when_ArraySlice_l166_233 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_233_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_233_2);
  assign _zz_when_ArraySlice_l166_233_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_233_3);
  assign _zz_when_ArraySlice_l166_233_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_233_3 = {2'd0, _zz_when_ArraySlice_l166_233_4};
  assign _zz__zz_when_ArraySlice_l112_233 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_233 = (_zz_when_ArraySlice_l113_233_1 - _zz_when_ArraySlice_l113_233_4);
  assign _zz_when_ArraySlice_l113_233_1 = (_zz_when_ArraySlice_l113_233_2 + _zz_when_ArraySlice_l113_233_3);
  assign _zz_when_ArraySlice_l113_233_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_233_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_233_4 = {1'd0, _zz_when_ArraySlice_l112_233};
  assign _zz__zz_when_ArraySlice_l173_233 = (_zz__zz_when_ArraySlice_l173_233_1 + _zz__zz_when_ArraySlice_l173_233_2);
  assign _zz__zz_when_ArraySlice_l173_233_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_233_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_233_3 = {1'd0, _zz_when_ArraySlice_l112_233};
  assign _zz_when_ArraySlice_l118_233_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_233 = _zz_when_ArraySlice_l118_233_1[5:0];
  assign _zz_when_ArraySlice_l173_233_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_233_1 = {1'd0, _zz_when_ArraySlice_l173_233_2};
  assign _zz_when_ArraySlice_l173_233_3 = (_zz_when_ArraySlice_l173_233_4 + _zz_when_ArraySlice_l173_233_9);
  assign _zz_when_ArraySlice_l173_233_4 = (_zz_when_ArraySlice_l173_233 - _zz_when_ArraySlice_l173_233_5);
  assign _zz_when_ArraySlice_l173_233_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_233_7);
  assign _zz_when_ArraySlice_l173_233_5 = {1'd0, _zz_when_ArraySlice_l173_233_6};
  assign _zz_when_ArraySlice_l173_233_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_233_7 = {2'd0, _zz_when_ArraySlice_l173_233_8};
  assign _zz_when_ArraySlice_l173_233_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_234 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_234_1);
  assign _zz_when_ArraySlice_l165_234_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_234_1 = {1'd0, _zz_when_ArraySlice_l165_234_2};
  assign _zz_when_ArraySlice_l166_234 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_234_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_234_2);
  assign _zz_when_ArraySlice_l166_234_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_234_3);
  assign _zz_when_ArraySlice_l166_234_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_234_3 = {1'd0, _zz_when_ArraySlice_l166_234_4};
  assign _zz__zz_when_ArraySlice_l112_234 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_234 = (_zz_when_ArraySlice_l113_234_1 - _zz_when_ArraySlice_l113_234_4);
  assign _zz_when_ArraySlice_l113_234_1 = (_zz_when_ArraySlice_l113_234_2 + _zz_when_ArraySlice_l113_234_3);
  assign _zz_when_ArraySlice_l113_234_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_234_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_234_4 = {1'd0, _zz_when_ArraySlice_l112_234};
  assign _zz__zz_when_ArraySlice_l173_234 = (_zz__zz_when_ArraySlice_l173_234_1 + _zz__zz_when_ArraySlice_l173_234_2);
  assign _zz__zz_when_ArraySlice_l173_234_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_234_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_234_3 = {1'd0, _zz_when_ArraySlice_l112_234};
  assign _zz_when_ArraySlice_l118_234_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_234 = _zz_when_ArraySlice_l118_234_1[5:0];
  assign _zz_when_ArraySlice_l173_234_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_234_1 = {1'd0, _zz_when_ArraySlice_l173_234_2};
  assign _zz_when_ArraySlice_l173_234_3 = (_zz_when_ArraySlice_l173_234_4 + _zz_when_ArraySlice_l173_234_9);
  assign _zz_when_ArraySlice_l173_234_4 = (_zz_when_ArraySlice_l173_234 - _zz_when_ArraySlice_l173_234_5);
  assign _zz_when_ArraySlice_l173_234_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_234_7);
  assign _zz_when_ArraySlice_l173_234_5 = {1'd0, _zz_when_ArraySlice_l173_234_6};
  assign _zz_when_ArraySlice_l173_234_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_234_7 = {1'd0, _zz_when_ArraySlice_l173_234_8};
  assign _zz_when_ArraySlice_l173_234_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_235 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_235_1);
  assign _zz_when_ArraySlice_l165_235_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_235_1 = {1'd0, _zz_when_ArraySlice_l165_235_2};
  assign _zz_when_ArraySlice_l166_235 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_235_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_235_2);
  assign _zz_when_ArraySlice_l166_235_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_235_3);
  assign _zz_when_ArraySlice_l166_235_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_235_3 = {1'd0, _zz_when_ArraySlice_l166_235_4};
  assign _zz__zz_when_ArraySlice_l112_235 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_235 = (_zz_when_ArraySlice_l113_235_1 - _zz_when_ArraySlice_l113_235_4);
  assign _zz_when_ArraySlice_l113_235_1 = (_zz_when_ArraySlice_l113_235_2 + _zz_when_ArraySlice_l113_235_3);
  assign _zz_when_ArraySlice_l113_235_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_235_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_235_4 = {1'd0, _zz_when_ArraySlice_l112_235};
  assign _zz__zz_when_ArraySlice_l173_235 = (_zz__zz_when_ArraySlice_l173_235_1 + _zz__zz_when_ArraySlice_l173_235_2);
  assign _zz__zz_when_ArraySlice_l173_235_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_235_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_235_3 = {1'd0, _zz_when_ArraySlice_l112_235};
  assign _zz_when_ArraySlice_l118_235_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_235 = _zz_when_ArraySlice_l118_235_1[5:0];
  assign _zz_when_ArraySlice_l173_235_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_235_1 = {1'd0, _zz_when_ArraySlice_l173_235_2};
  assign _zz_when_ArraySlice_l173_235_3 = (_zz_when_ArraySlice_l173_235_4 + _zz_when_ArraySlice_l173_235_9);
  assign _zz_when_ArraySlice_l173_235_4 = (_zz_when_ArraySlice_l173_235 - _zz_when_ArraySlice_l173_235_5);
  assign _zz_when_ArraySlice_l173_235_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_235_7);
  assign _zz_when_ArraySlice_l173_235_5 = {1'd0, _zz_when_ArraySlice_l173_235_6};
  assign _zz_when_ArraySlice_l173_235_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_235_7 = {1'd0, _zz_when_ArraySlice_l173_235_8};
  assign _zz_when_ArraySlice_l173_235_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_236 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_236_1);
  assign _zz_when_ArraySlice_l165_236_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_236 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_236_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_236_2);
  assign _zz_when_ArraySlice_l166_236_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_236_3);
  assign _zz_when_ArraySlice_l166_236_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_236 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_236 = (_zz_when_ArraySlice_l113_236_1 - _zz_when_ArraySlice_l113_236_4);
  assign _zz_when_ArraySlice_l113_236_1 = (_zz_when_ArraySlice_l113_236_2 + _zz_when_ArraySlice_l113_236_3);
  assign _zz_when_ArraySlice_l113_236_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_236_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_236_4 = {1'd0, _zz_when_ArraySlice_l112_236};
  assign _zz__zz_when_ArraySlice_l173_236 = (_zz__zz_when_ArraySlice_l173_236_1 + _zz__zz_when_ArraySlice_l173_236_2);
  assign _zz__zz_when_ArraySlice_l173_236_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_236_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_236_3 = {1'd0, _zz_when_ArraySlice_l112_236};
  assign _zz_when_ArraySlice_l118_236_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_236 = _zz_when_ArraySlice_l118_236_1[5:0];
  assign _zz_when_ArraySlice_l173_236_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_236_1 = {1'd0, _zz_when_ArraySlice_l173_236_2};
  assign _zz_when_ArraySlice_l173_236_3 = (_zz_when_ArraySlice_l173_236_4 + _zz_when_ArraySlice_l173_236_8);
  assign _zz_when_ArraySlice_l173_236_4 = (_zz_when_ArraySlice_l173_236 - _zz_when_ArraySlice_l173_236_5);
  assign _zz_when_ArraySlice_l173_236_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_236_7);
  assign _zz_when_ArraySlice_l173_236_5 = {1'd0, _zz_when_ArraySlice_l173_236_6};
  assign _zz_when_ArraySlice_l173_236_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_236_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_237 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_237_1);
  assign _zz_when_ArraySlice_l165_237_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_237_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_237 = {1'd0, _zz_when_ArraySlice_l166_237_1};
  assign _zz_when_ArraySlice_l166_237_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_237_3);
  assign _zz_when_ArraySlice_l166_237_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_237_4);
  assign _zz_when_ArraySlice_l166_237_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_237 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_237 = (_zz_when_ArraySlice_l113_237_1 - _zz_when_ArraySlice_l113_237_4);
  assign _zz_when_ArraySlice_l113_237_1 = (_zz_when_ArraySlice_l113_237_2 + _zz_when_ArraySlice_l113_237_3);
  assign _zz_when_ArraySlice_l113_237_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_237_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_237_4 = {1'd0, _zz_when_ArraySlice_l112_237};
  assign _zz__zz_when_ArraySlice_l173_237 = (_zz__zz_when_ArraySlice_l173_237_1 + _zz__zz_when_ArraySlice_l173_237_2);
  assign _zz__zz_when_ArraySlice_l173_237_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_237_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_237_3 = {1'd0, _zz_when_ArraySlice_l112_237};
  assign _zz_when_ArraySlice_l118_237_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_237 = _zz_when_ArraySlice_l118_237_1[5:0];
  assign _zz_when_ArraySlice_l173_237_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_237_1 = {2'd0, _zz_when_ArraySlice_l173_237_2};
  assign _zz_when_ArraySlice_l173_237_3 = (_zz_when_ArraySlice_l173_237_4 + _zz_when_ArraySlice_l173_237_8);
  assign _zz_when_ArraySlice_l173_237_4 = (_zz_when_ArraySlice_l173_237 - _zz_when_ArraySlice_l173_237_5);
  assign _zz_when_ArraySlice_l173_237_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_237_7);
  assign _zz_when_ArraySlice_l173_237_5 = {1'd0, _zz_when_ArraySlice_l173_237_6};
  assign _zz_when_ArraySlice_l173_237_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_237_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_238 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_238_1);
  assign _zz_when_ArraySlice_l165_238_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_238_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_238 = {1'd0, _zz_when_ArraySlice_l166_238_1};
  assign _zz_when_ArraySlice_l166_238_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_238_3);
  assign _zz_when_ArraySlice_l166_238_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_238_4);
  assign _zz_when_ArraySlice_l166_238_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_238 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_238 = (_zz_when_ArraySlice_l113_238_1 - _zz_when_ArraySlice_l113_238_4);
  assign _zz_when_ArraySlice_l113_238_1 = (_zz_when_ArraySlice_l113_238_2 + _zz_when_ArraySlice_l113_238_3);
  assign _zz_when_ArraySlice_l113_238_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_238_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_238_4 = {1'd0, _zz_when_ArraySlice_l112_238};
  assign _zz__zz_when_ArraySlice_l173_238 = (_zz__zz_when_ArraySlice_l173_238_1 + _zz__zz_when_ArraySlice_l173_238_2);
  assign _zz__zz_when_ArraySlice_l173_238_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_238_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_238_3 = {1'd0, _zz_when_ArraySlice_l112_238};
  assign _zz_when_ArraySlice_l118_238_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_238 = _zz_when_ArraySlice_l118_238_1[5:0];
  assign _zz_when_ArraySlice_l173_238_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_238_1 = {2'd0, _zz_when_ArraySlice_l173_238_2};
  assign _zz_when_ArraySlice_l173_238_3 = (_zz_when_ArraySlice_l173_238_4 + _zz_when_ArraySlice_l173_238_8);
  assign _zz_when_ArraySlice_l173_238_4 = (_zz_when_ArraySlice_l173_238 - _zz_when_ArraySlice_l173_238_5);
  assign _zz_when_ArraySlice_l173_238_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_238_7);
  assign _zz_when_ArraySlice_l173_238_5 = {1'd0, _zz_when_ArraySlice_l173_238_6};
  assign _zz_when_ArraySlice_l173_238_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_238_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_239 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_239_1);
  assign _zz_when_ArraySlice_l165_239_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_239_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_239 = {2'd0, _zz_when_ArraySlice_l166_239_1};
  assign _zz_when_ArraySlice_l166_239_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_239_3);
  assign _zz_when_ArraySlice_l166_239_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_239_4);
  assign _zz_when_ArraySlice_l166_239_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_239 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_239 = (_zz_when_ArraySlice_l113_239_1 - _zz_when_ArraySlice_l113_239_4);
  assign _zz_when_ArraySlice_l113_239_1 = (_zz_when_ArraySlice_l113_239_2 + _zz_when_ArraySlice_l113_239_3);
  assign _zz_when_ArraySlice_l113_239_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_239_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_239_4 = {1'd0, _zz_when_ArraySlice_l112_239};
  assign _zz__zz_when_ArraySlice_l173_239 = (_zz__zz_when_ArraySlice_l173_239_1 + _zz__zz_when_ArraySlice_l173_239_2);
  assign _zz__zz_when_ArraySlice_l173_239_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_239_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_239_3 = {1'd0, _zz_when_ArraySlice_l112_239};
  assign _zz_when_ArraySlice_l118_239_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_239 = _zz_when_ArraySlice_l118_239_1[5:0];
  assign _zz_when_ArraySlice_l173_239_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_239_1 = {3'd0, _zz_when_ArraySlice_l173_239_2};
  assign _zz_when_ArraySlice_l173_239_3 = (_zz_when_ArraySlice_l173_239_4 + _zz_when_ArraySlice_l173_239_8);
  assign _zz_when_ArraySlice_l173_239_4 = (_zz_when_ArraySlice_l173_239 - _zz_when_ArraySlice_l173_239_5);
  assign _zz_when_ArraySlice_l173_239_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_239_7);
  assign _zz_when_ArraySlice_l173_239_5 = {1'd0, _zz_when_ArraySlice_l173_239_6};
  assign _zz_when_ArraySlice_l173_239_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_239_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l268_1_1 = (_zz_when_ArraySlice_l268_1_2 + _zz_when_ArraySlice_l268_1_7);
  assign _zz_when_ArraySlice_l268_1_2 = (_zz_when_ArraySlice_l268_1_3 + _zz_when_ArraySlice_l268_1_5);
  assign _zz_when_ArraySlice_l268_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l268_1_4);
  assign _zz_when_ArraySlice_l268_1_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l268_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l268_1_5 = {5'd0, _zz_when_ArraySlice_l268_1_6};
  assign _zz_when_ArraySlice_l268_1_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l268_1_7 = {2'd0, _zz_when_ArraySlice_l268_1_8};
  assign _zz_selectReadFifo_1_47 = 1'b1;
  assign _zz_selectReadFifo_1_46 = {5'd0, _zz_selectReadFifo_1_47};
  assign _zz_when_ArraySlice_l272_1_1 = (_zz_when_ArraySlice_l272_1_2 % aReg);
  assign _zz_when_ArraySlice_l272_1_2 = (handshakeTimes_1_value + _zz_when_ArraySlice_l272_1_3);
  assign _zz_when_ArraySlice_l272_1_4 = 1'b1;
  assign _zz_when_ArraySlice_l272_1_3 = {12'd0, _zz_when_ArraySlice_l272_1_4};
  assign _zz_when_ArraySlice_l276_1_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l276_1_3);
  assign _zz_when_ArraySlice_l276_1_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l276_1_3 = {2'd0, _zz_when_ArraySlice_l276_1_4};
  assign _zz_when_ArraySlice_l277_1_2 = (_zz_when_ArraySlice_l277_1_3 - _zz_when_ArraySlice_l277_1_4);
  assign _zz_when_ArraySlice_l277_1_1 = {7'd0, _zz_when_ArraySlice_l277_1_2};
  assign _zz_when_ArraySlice_l277_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l277_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l277_1_4 = {5'd0, _zz_when_ArraySlice_l277_1_5};
  assign _zz__zz_when_ArraySlice_l94_28 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_28 = (_zz_when_ArraySlice_l95_28_1 - _zz_when_ArraySlice_l95_28_4);
  assign _zz_when_ArraySlice_l95_28_1 = (_zz_when_ArraySlice_l95_28_2 + _zz_when_ArraySlice_l95_28_3);
  assign _zz_when_ArraySlice_l95_28_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_28_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_28_4 = {1'd0, _zz_when_ArraySlice_l94_28};
  assign _zz__zz_when_ArraySlice_l279_1_1 = (_zz__zz_when_ArraySlice_l279_1_2 + _zz__zz_when_ArraySlice_l279_1_3);
  assign _zz__zz_when_ArraySlice_l279_1_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l279_1_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l279_1_4 = {1'd0, _zz_when_ArraySlice_l94_28};
  assign _zz_when_ArraySlice_l99_28_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_28 = _zz_when_ArraySlice_l99_28_1[5:0];
  assign _zz_when_ArraySlice_l279_1_1 = (outSliceNumb_1_value + _zz_when_ArraySlice_l279_1_2);
  assign _zz_when_ArraySlice_l279_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l279_1_2 = {6'd0, _zz_when_ArraySlice_l279_1_3};
  assign _zz_when_ArraySlice_l279_1_4 = (_zz_when_ArraySlice_l279_1 / aReg);
  assign _zz_selectReadFifo_1_48 = (selectReadFifo_1 - _zz_selectReadFifo_1_49);
  assign _zz_selectReadFifo_1_49 = {3'd0, bReg};
  assign _zz_selectReadFifo_1_51 = 1'b1;
  assign _zz_selectReadFifo_1_50 = {5'd0, _zz_selectReadFifo_1_51};
  assign _zz_selectReadFifo_1_52 = (selectReadFifo_1 + _zz_selectReadFifo_1_53);
  assign _zz_selectReadFifo_1_53 = (3'b111 * bReg);
  assign _zz_selectReadFifo_1_55 = 1'b1;
  assign _zz_selectReadFifo_1_54 = {5'd0, _zz_selectReadFifo_1_55};
  assign _zz_when_ArraySlice_l165_240 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_240_1);
  assign _zz_when_ArraySlice_l165_240_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_240_1 = {3'd0, _zz_when_ArraySlice_l165_240_2};
  assign _zz_when_ArraySlice_l166_240 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_240_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_240_3);
  assign _zz_when_ArraySlice_l166_240_1 = {1'd0, _zz_when_ArraySlice_l166_240_2};
  assign _zz_when_ArraySlice_l166_240_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_240_4);
  assign _zz_when_ArraySlice_l166_240_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_240_4 = {3'd0, _zz_when_ArraySlice_l166_240_5};
  assign _zz__zz_when_ArraySlice_l112_240 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_240 = (_zz_when_ArraySlice_l113_240_1 - _zz_when_ArraySlice_l113_240_4);
  assign _zz_when_ArraySlice_l113_240_1 = (_zz_when_ArraySlice_l113_240_2 + _zz_when_ArraySlice_l113_240_3);
  assign _zz_when_ArraySlice_l113_240_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_240_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_240_4 = {1'd0, _zz_when_ArraySlice_l112_240};
  assign _zz__zz_when_ArraySlice_l173_240 = (_zz__zz_when_ArraySlice_l173_240_1 + _zz__zz_when_ArraySlice_l173_240_2);
  assign _zz__zz_when_ArraySlice_l173_240_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_240_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_240_3 = {1'd0, _zz_when_ArraySlice_l112_240};
  assign _zz_when_ArraySlice_l118_240_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_240 = _zz_when_ArraySlice_l118_240_1[5:0];
  assign _zz_when_ArraySlice_l173_240_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_240_2 = (_zz_when_ArraySlice_l173_240_3 + _zz_when_ArraySlice_l173_240_8);
  assign _zz_when_ArraySlice_l173_240_3 = (_zz_when_ArraySlice_l173_240 - _zz_when_ArraySlice_l173_240_4);
  assign _zz_when_ArraySlice_l173_240_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_240_6);
  assign _zz_when_ArraySlice_l173_240_4 = {1'd0, _zz_when_ArraySlice_l173_240_5};
  assign _zz_when_ArraySlice_l173_240_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_240_6 = {3'd0, _zz_when_ArraySlice_l173_240_7};
  assign _zz_when_ArraySlice_l173_240_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_241 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_241_1);
  assign _zz_when_ArraySlice_l165_241_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_241_1 = {2'd0, _zz_when_ArraySlice_l165_241_2};
  assign _zz_when_ArraySlice_l166_241 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_241_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_241_2);
  assign _zz_when_ArraySlice_l166_241_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_241_3);
  assign _zz_when_ArraySlice_l166_241_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_241_3 = {2'd0, _zz_when_ArraySlice_l166_241_4};
  assign _zz__zz_when_ArraySlice_l112_241 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_241 = (_zz_when_ArraySlice_l113_241_1 - _zz_when_ArraySlice_l113_241_4);
  assign _zz_when_ArraySlice_l113_241_1 = (_zz_when_ArraySlice_l113_241_2 + _zz_when_ArraySlice_l113_241_3);
  assign _zz_when_ArraySlice_l113_241_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_241_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_241_4 = {1'd0, _zz_when_ArraySlice_l112_241};
  assign _zz__zz_when_ArraySlice_l173_241 = (_zz__zz_when_ArraySlice_l173_241_1 + _zz__zz_when_ArraySlice_l173_241_2);
  assign _zz__zz_when_ArraySlice_l173_241_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_241_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_241_3 = {1'd0, _zz_when_ArraySlice_l112_241};
  assign _zz_when_ArraySlice_l118_241_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_241 = _zz_when_ArraySlice_l118_241_1[5:0];
  assign _zz_when_ArraySlice_l173_241_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_241_1 = {1'd0, _zz_when_ArraySlice_l173_241_2};
  assign _zz_when_ArraySlice_l173_241_3 = (_zz_when_ArraySlice_l173_241_4 + _zz_when_ArraySlice_l173_241_9);
  assign _zz_when_ArraySlice_l173_241_4 = (_zz_when_ArraySlice_l173_241 - _zz_when_ArraySlice_l173_241_5);
  assign _zz_when_ArraySlice_l173_241_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_241_7);
  assign _zz_when_ArraySlice_l173_241_5 = {1'd0, _zz_when_ArraySlice_l173_241_6};
  assign _zz_when_ArraySlice_l173_241_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_241_7 = {2'd0, _zz_when_ArraySlice_l173_241_8};
  assign _zz_when_ArraySlice_l173_241_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_242 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_242_1);
  assign _zz_when_ArraySlice_l165_242_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_242_1 = {1'd0, _zz_when_ArraySlice_l165_242_2};
  assign _zz_when_ArraySlice_l166_242 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_242_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_242_2);
  assign _zz_when_ArraySlice_l166_242_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_242_3);
  assign _zz_when_ArraySlice_l166_242_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_242_3 = {1'd0, _zz_when_ArraySlice_l166_242_4};
  assign _zz__zz_when_ArraySlice_l112_242 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_242 = (_zz_when_ArraySlice_l113_242_1 - _zz_when_ArraySlice_l113_242_4);
  assign _zz_when_ArraySlice_l113_242_1 = (_zz_when_ArraySlice_l113_242_2 + _zz_when_ArraySlice_l113_242_3);
  assign _zz_when_ArraySlice_l113_242_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_242_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_242_4 = {1'd0, _zz_when_ArraySlice_l112_242};
  assign _zz__zz_when_ArraySlice_l173_242 = (_zz__zz_when_ArraySlice_l173_242_1 + _zz__zz_when_ArraySlice_l173_242_2);
  assign _zz__zz_when_ArraySlice_l173_242_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_242_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_242_3 = {1'd0, _zz_when_ArraySlice_l112_242};
  assign _zz_when_ArraySlice_l118_242_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_242 = _zz_when_ArraySlice_l118_242_1[5:0];
  assign _zz_when_ArraySlice_l173_242_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_242_1 = {1'd0, _zz_when_ArraySlice_l173_242_2};
  assign _zz_when_ArraySlice_l173_242_3 = (_zz_when_ArraySlice_l173_242_4 + _zz_when_ArraySlice_l173_242_9);
  assign _zz_when_ArraySlice_l173_242_4 = (_zz_when_ArraySlice_l173_242 - _zz_when_ArraySlice_l173_242_5);
  assign _zz_when_ArraySlice_l173_242_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_242_7);
  assign _zz_when_ArraySlice_l173_242_5 = {1'd0, _zz_when_ArraySlice_l173_242_6};
  assign _zz_when_ArraySlice_l173_242_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_242_7 = {1'd0, _zz_when_ArraySlice_l173_242_8};
  assign _zz_when_ArraySlice_l173_242_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_243 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_243_1);
  assign _zz_when_ArraySlice_l165_243_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_243_1 = {1'd0, _zz_when_ArraySlice_l165_243_2};
  assign _zz_when_ArraySlice_l166_243 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_243_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_243_2);
  assign _zz_when_ArraySlice_l166_243_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_243_3);
  assign _zz_when_ArraySlice_l166_243_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_243_3 = {1'd0, _zz_when_ArraySlice_l166_243_4};
  assign _zz__zz_when_ArraySlice_l112_243 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_243 = (_zz_when_ArraySlice_l113_243_1 - _zz_when_ArraySlice_l113_243_4);
  assign _zz_when_ArraySlice_l113_243_1 = (_zz_when_ArraySlice_l113_243_2 + _zz_when_ArraySlice_l113_243_3);
  assign _zz_when_ArraySlice_l113_243_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_243_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_243_4 = {1'd0, _zz_when_ArraySlice_l112_243};
  assign _zz__zz_when_ArraySlice_l173_243 = (_zz__zz_when_ArraySlice_l173_243_1 + _zz__zz_when_ArraySlice_l173_243_2);
  assign _zz__zz_when_ArraySlice_l173_243_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_243_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_243_3 = {1'd0, _zz_when_ArraySlice_l112_243};
  assign _zz_when_ArraySlice_l118_243_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_243 = _zz_when_ArraySlice_l118_243_1[5:0];
  assign _zz_when_ArraySlice_l173_243_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_243_1 = {1'd0, _zz_when_ArraySlice_l173_243_2};
  assign _zz_when_ArraySlice_l173_243_3 = (_zz_when_ArraySlice_l173_243_4 + _zz_when_ArraySlice_l173_243_9);
  assign _zz_when_ArraySlice_l173_243_4 = (_zz_when_ArraySlice_l173_243 - _zz_when_ArraySlice_l173_243_5);
  assign _zz_when_ArraySlice_l173_243_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_243_7);
  assign _zz_when_ArraySlice_l173_243_5 = {1'd0, _zz_when_ArraySlice_l173_243_6};
  assign _zz_when_ArraySlice_l173_243_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_243_7 = {1'd0, _zz_when_ArraySlice_l173_243_8};
  assign _zz_when_ArraySlice_l173_243_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_244 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_244_1);
  assign _zz_when_ArraySlice_l165_244_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_244 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_244_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_244_2);
  assign _zz_when_ArraySlice_l166_244_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_244_3);
  assign _zz_when_ArraySlice_l166_244_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_244 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_244 = (_zz_when_ArraySlice_l113_244_1 - _zz_when_ArraySlice_l113_244_4);
  assign _zz_when_ArraySlice_l113_244_1 = (_zz_when_ArraySlice_l113_244_2 + _zz_when_ArraySlice_l113_244_3);
  assign _zz_when_ArraySlice_l113_244_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_244_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_244_4 = {1'd0, _zz_when_ArraySlice_l112_244};
  assign _zz__zz_when_ArraySlice_l173_244 = (_zz__zz_when_ArraySlice_l173_244_1 + _zz__zz_when_ArraySlice_l173_244_2);
  assign _zz__zz_when_ArraySlice_l173_244_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_244_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_244_3 = {1'd0, _zz_when_ArraySlice_l112_244};
  assign _zz_when_ArraySlice_l118_244_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_244 = _zz_when_ArraySlice_l118_244_1[5:0];
  assign _zz_when_ArraySlice_l173_244_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_244_1 = {1'd0, _zz_when_ArraySlice_l173_244_2};
  assign _zz_when_ArraySlice_l173_244_3 = (_zz_when_ArraySlice_l173_244_4 + _zz_when_ArraySlice_l173_244_8);
  assign _zz_when_ArraySlice_l173_244_4 = (_zz_when_ArraySlice_l173_244 - _zz_when_ArraySlice_l173_244_5);
  assign _zz_when_ArraySlice_l173_244_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_244_7);
  assign _zz_when_ArraySlice_l173_244_5 = {1'd0, _zz_when_ArraySlice_l173_244_6};
  assign _zz_when_ArraySlice_l173_244_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_244_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_245 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_245_1);
  assign _zz_when_ArraySlice_l165_245_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_245_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_245 = {1'd0, _zz_when_ArraySlice_l166_245_1};
  assign _zz_when_ArraySlice_l166_245_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_245_3);
  assign _zz_when_ArraySlice_l166_245_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_245_4);
  assign _zz_when_ArraySlice_l166_245_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_245 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_245 = (_zz_when_ArraySlice_l113_245_1 - _zz_when_ArraySlice_l113_245_4);
  assign _zz_when_ArraySlice_l113_245_1 = (_zz_when_ArraySlice_l113_245_2 + _zz_when_ArraySlice_l113_245_3);
  assign _zz_when_ArraySlice_l113_245_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_245_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_245_4 = {1'd0, _zz_when_ArraySlice_l112_245};
  assign _zz__zz_when_ArraySlice_l173_245 = (_zz__zz_when_ArraySlice_l173_245_1 + _zz__zz_when_ArraySlice_l173_245_2);
  assign _zz__zz_when_ArraySlice_l173_245_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_245_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_245_3 = {1'd0, _zz_when_ArraySlice_l112_245};
  assign _zz_when_ArraySlice_l118_245_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_245 = _zz_when_ArraySlice_l118_245_1[5:0];
  assign _zz_when_ArraySlice_l173_245_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_245_1 = {2'd0, _zz_when_ArraySlice_l173_245_2};
  assign _zz_when_ArraySlice_l173_245_3 = (_zz_when_ArraySlice_l173_245_4 + _zz_when_ArraySlice_l173_245_8);
  assign _zz_when_ArraySlice_l173_245_4 = (_zz_when_ArraySlice_l173_245 - _zz_when_ArraySlice_l173_245_5);
  assign _zz_when_ArraySlice_l173_245_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_245_7);
  assign _zz_when_ArraySlice_l173_245_5 = {1'd0, _zz_when_ArraySlice_l173_245_6};
  assign _zz_when_ArraySlice_l173_245_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_245_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_246 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_246_1);
  assign _zz_when_ArraySlice_l165_246_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_246_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_246 = {1'd0, _zz_when_ArraySlice_l166_246_1};
  assign _zz_when_ArraySlice_l166_246_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_246_3);
  assign _zz_when_ArraySlice_l166_246_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_246_4);
  assign _zz_when_ArraySlice_l166_246_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_246 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_246 = (_zz_when_ArraySlice_l113_246_1 - _zz_when_ArraySlice_l113_246_4);
  assign _zz_when_ArraySlice_l113_246_1 = (_zz_when_ArraySlice_l113_246_2 + _zz_when_ArraySlice_l113_246_3);
  assign _zz_when_ArraySlice_l113_246_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_246_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_246_4 = {1'd0, _zz_when_ArraySlice_l112_246};
  assign _zz__zz_when_ArraySlice_l173_246 = (_zz__zz_when_ArraySlice_l173_246_1 + _zz__zz_when_ArraySlice_l173_246_2);
  assign _zz__zz_when_ArraySlice_l173_246_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_246_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_246_3 = {1'd0, _zz_when_ArraySlice_l112_246};
  assign _zz_when_ArraySlice_l118_246_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_246 = _zz_when_ArraySlice_l118_246_1[5:0];
  assign _zz_when_ArraySlice_l173_246_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_246_1 = {2'd0, _zz_when_ArraySlice_l173_246_2};
  assign _zz_when_ArraySlice_l173_246_3 = (_zz_when_ArraySlice_l173_246_4 + _zz_when_ArraySlice_l173_246_8);
  assign _zz_when_ArraySlice_l173_246_4 = (_zz_when_ArraySlice_l173_246 - _zz_when_ArraySlice_l173_246_5);
  assign _zz_when_ArraySlice_l173_246_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_246_7);
  assign _zz_when_ArraySlice_l173_246_5 = {1'd0, _zz_when_ArraySlice_l173_246_6};
  assign _zz_when_ArraySlice_l173_246_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_246_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_247 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_247_1);
  assign _zz_when_ArraySlice_l165_247_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_247_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_247 = {2'd0, _zz_when_ArraySlice_l166_247_1};
  assign _zz_when_ArraySlice_l166_247_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_247_3);
  assign _zz_when_ArraySlice_l166_247_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_247_4);
  assign _zz_when_ArraySlice_l166_247_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_247 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_247 = (_zz_when_ArraySlice_l113_247_1 - _zz_when_ArraySlice_l113_247_4);
  assign _zz_when_ArraySlice_l113_247_1 = (_zz_when_ArraySlice_l113_247_2 + _zz_when_ArraySlice_l113_247_3);
  assign _zz_when_ArraySlice_l113_247_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_247_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_247_4 = {1'd0, _zz_when_ArraySlice_l112_247};
  assign _zz__zz_when_ArraySlice_l173_247 = (_zz__zz_when_ArraySlice_l173_247_1 + _zz__zz_when_ArraySlice_l173_247_2);
  assign _zz__zz_when_ArraySlice_l173_247_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_247_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_247_3 = {1'd0, _zz_when_ArraySlice_l112_247};
  assign _zz_when_ArraySlice_l118_247_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_247 = _zz_when_ArraySlice_l118_247_1[5:0];
  assign _zz_when_ArraySlice_l173_247_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_247_1 = {3'd0, _zz_when_ArraySlice_l173_247_2};
  assign _zz_when_ArraySlice_l173_247_3 = (_zz_when_ArraySlice_l173_247_4 + _zz_when_ArraySlice_l173_247_8);
  assign _zz_when_ArraySlice_l173_247_4 = (_zz_when_ArraySlice_l173_247 - _zz_when_ArraySlice_l173_247_5);
  assign _zz_when_ArraySlice_l173_247_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_247_7);
  assign _zz_when_ArraySlice_l173_247_5 = {1'd0, _zz_when_ArraySlice_l173_247_6};
  assign _zz_when_ArraySlice_l173_247_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_247_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l288_1_1 = (_zz_when_ArraySlice_l288_1_2 + _zz_when_ArraySlice_l288_1_7);
  assign _zz_when_ArraySlice_l288_1_2 = (_zz_when_ArraySlice_l288_1_3 + _zz_when_ArraySlice_l288_1_5);
  assign _zz_when_ArraySlice_l288_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l288_1_4);
  assign _zz_when_ArraySlice_l288_1_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l288_1_5 = {5'd0, _zz_when_ArraySlice_l288_1_6};
  assign _zz_when_ArraySlice_l288_1_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l288_1_7 = {2'd0, _zz_when_ArraySlice_l288_1_8};
  assign _zz_selectReadFifo_1_57 = 1'b1;
  assign _zz_selectReadFifo_1_56 = {5'd0, _zz_selectReadFifo_1_57};
  assign _zz_when_ArraySlice_l292_1_1 = (_zz_when_ArraySlice_l292_1_2 % aReg);
  assign _zz_when_ArraySlice_l292_1_2 = (handshakeTimes_1_value + _zz_when_ArraySlice_l292_1_3);
  assign _zz_when_ArraySlice_l292_1_4 = 1'b1;
  assign _zz_when_ArraySlice_l292_1_3 = {12'd0, _zz_when_ArraySlice_l292_1_4};
  assign _zz_when_ArraySlice_l303_1_2 = (_zz_when_ArraySlice_l303_1_3 - _zz_when_ArraySlice_l303_1_4);
  assign _zz_when_ArraySlice_l303_1_1 = {7'd0, _zz_when_ArraySlice_l303_1_2};
  assign _zz_when_ArraySlice_l303_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l303_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l303_1_4 = {5'd0, _zz_when_ArraySlice_l303_1_5};
  assign _zz__zz_when_ArraySlice_l94_29 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_29 = (_zz_when_ArraySlice_l95_29_1 - _zz_when_ArraySlice_l95_29_4);
  assign _zz_when_ArraySlice_l95_29_1 = (_zz_when_ArraySlice_l95_29_2 + _zz_when_ArraySlice_l95_29_3);
  assign _zz_when_ArraySlice_l95_29_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_29_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_29_4 = {1'd0, _zz_when_ArraySlice_l94_29};
  assign _zz__zz_when_ArraySlice_l304_1_1 = (_zz__zz_when_ArraySlice_l304_1_2 + _zz__zz_when_ArraySlice_l304_1_3);
  assign _zz__zz_when_ArraySlice_l304_1_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l304_1_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l304_1_4 = {1'd0, _zz_when_ArraySlice_l94_29};
  assign _zz_when_ArraySlice_l99_29_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_29 = _zz_when_ArraySlice_l99_29_1[5:0];
  assign _zz_when_ArraySlice_l304_1_1 = (outSliceNumb_1_value + _zz_when_ArraySlice_l304_1_2);
  assign _zz_when_ArraySlice_l304_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l304_1_2 = {6'd0, _zz_when_ArraySlice_l304_1_3};
  assign _zz_when_ArraySlice_l304_1_4 = (_zz_when_ArraySlice_l304_1 / aReg);
  assign _zz_selectReadFifo_1_58 = (selectReadFifo_1 - _zz_selectReadFifo_1_59);
  assign _zz_selectReadFifo_1_59 = {3'd0, bReg};
  assign _zz_selectReadFifo_1_61 = 1'b1;
  assign _zz_selectReadFifo_1_60 = {5'd0, _zz_selectReadFifo_1_61};
  assign _zz_when_ArraySlice_l165_248 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_248_1);
  assign _zz_when_ArraySlice_l165_248_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_248_1 = {3'd0, _zz_when_ArraySlice_l165_248_2};
  assign _zz_when_ArraySlice_l166_248 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_248_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_248_3);
  assign _zz_when_ArraySlice_l166_248_1 = {1'd0, _zz_when_ArraySlice_l166_248_2};
  assign _zz_when_ArraySlice_l166_248_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_248_4);
  assign _zz_when_ArraySlice_l166_248_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_248_4 = {3'd0, _zz_when_ArraySlice_l166_248_5};
  assign _zz__zz_when_ArraySlice_l112_248 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_248 = (_zz_when_ArraySlice_l113_248_1 - _zz_when_ArraySlice_l113_248_4);
  assign _zz_when_ArraySlice_l113_248_1 = (_zz_when_ArraySlice_l113_248_2 + _zz_when_ArraySlice_l113_248_3);
  assign _zz_when_ArraySlice_l113_248_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_248_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_248_4 = {1'd0, _zz_when_ArraySlice_l112_248};
  assign _zz__zz_when_ArraySlice_l173_248 = (_zz__zz_when_ArraySlice_l173_248_1 + _zz__zz_when_ArraySlice_l173_248_2);
  assign _zz__zz_when_ArraySlice_l173_248_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_248_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_248_3 = {1'd0, _zz_when_ArraySlice_l112_248};
  assign _zz_when_ArraySlice_l118_248_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_248 = _zz_when_ArraySlice_l118_248_1[5:0];
  assign _zz_when_ArraySlice_l173_248_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_248_2 = (_zz_when_ArraySlice_l173_248_3 + _zz_when_ArraySlice_l173_248_8);
  assign _zz_when_ArraySlice_l173_248_3 = (_zz_when_ArraySlice_l173_248 - _zz_when_ArraySlice_l173_248_4);
  assign _zz_when_ArraySlice_l173_248_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_248_6);
  assign _zz_when_ArraySlice_l173_248_4 = {1'd0, _zz_when_ArraySlice_l173_248_5};
  assign _zz_when_ArraySlice_l173_248_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_248_6 = {3'd0, _zz_when_ArraySlice_l173_248_7};
  assign _zz_when_ArraySlice_l173_248_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_249 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_249_1);
  assign _zz_when_ArraySlice_l165_249_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_249_1 = {2'd0, _zz_when_ArraySlice_l165_249_2};
  assign _zz_when_ArraySlice_l166_249 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_249_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_249_2);
  assign _zz_when_ArraySlice_l166_249_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_249_3);
  assign _zz_when_ArraySlice_l166_249_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_249_3 = {2'd0, _zz_when_ArraySlice_l166_249_4};
  assign _zz__zz_when_ArraySlice_l112_249 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_249 = (_zz_when_ArraySlice_l113_249_1 - _zz_when_ArraySlice_l113_249_4);
  assign _zz_when_ArraySlice_l113_249_1 = (_zz_when_ArraySlice_l113_249_2 + _zz_when_ArraySlice_l113_249_3);
  assign _zz_when_ArraySlice_l113_249_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_249_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_249_4 = {1'd0, _zz_when_ArraySlice_l112_249};
  assign _zz__zz_when_ArraySlice_l173_249 = (_zz__zz_when_ArraySlice_l173_249_1 + _zz__zz_when_ArraySlice_l173_249_2);
  assign _zz__zz_when_ArraySlice_l173_249_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_249_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_249_3 = {1'd0, _zz_when_ArraySlice_l112_249};
  assign _zz_when_ArraySlice_l118_249_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_249 = _zz_when_ArraySlice_l118_249_1[5:0];
  assign _zz_when_ArraySlice_l173_249_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_249_1 = {1'd0, _zz_when_ArraySlice_l173_249_2};
  assign _zz_when_ArraySlice_l173_249_3 = (_zz_when_ArraySlice_l173_249_4 + _zz_when_ArraySlice_l173_249_9);
  assign _zz_when_ArraySlice_l173_249_4 = (_zz_when_ArraySlice_l173_249 - _zz_when_ArraySlice_l173_249_5);
  assign _zz_when_ArraySlice_l173_249_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_249_7);
  assign _zz_when_ArraySlice_l173_249_5 = {1'd0, _zz_when_ArraySlice_l173_249_6};
  assign _zz_when_ArraySlice_l173_249_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_249_7 = {2'd0, _zz_when_ArraySlice_l173_249_8};
  assign _zz_when_ArraySlice_l173_249_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_250 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_250_1);
  assign _zz_when_ArraySlice_l165_250_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_250_1 = {1'd0, _zz_when_ArraySlice_l165_250_2};
  assign _zz_when_ArraySlice_l166_250 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_250_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_250_2);
  assign _zz_when_ArraySlice_l166_250_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_250_3);
  assign _zz_when_ArraySlice_l166_250_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_250_3 = {1'd0, _zz_when_ArraySlice_l166_250_4};
  assign _zz__zz_when_ArraySlice_l112_250 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_250 = (_zz_when_ArraySlice_l113_250_1 - _zz_when_ArraySlice_l113_250_4);
  assign _zz_when_ArraySlice_l113_250_1 = (_zz_when_ArraySlice_l113_250_2 + _zz_when_ArraySlice_l113_250_3);
  assign _zz_when_ArraySlice_l113_250_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_250_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_250_4 = {1'd0, _zz_when_ArraySlice_l112_250};
  assign _zz__zz_when_ArraySlice_l173_250 = (_zz__zz_when_ArraySlice_l173_250_1 + _zz__zz_when_ArraySlice_l173_250_2);
  assign _zz__zz_when_ArraySlice_l173_250_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_250_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_250_3 = {1'd0, _zz_when_ArraySlice_l112_250};
  assign _zz_when_ArraySlice_l118_250_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_250 = _zz_when_ArraySlice_l118_250_1[5:0];
  assign _zz_when_ArraySlice_l173_250_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_250_1 = {1'd0, _zz_when_ArraySlice_l173_250_2};
  assign _zz_when_ArraySlice_l173_250_3 = (_zz_when_ArraySlice_l173_250_4 + _zz_when_ArraySlice_l173_250_9);
  assign _zz_when_ArraySlice_l173_250_4 = (_zz_when_ArraySlice_l173_250 - _zz_when_ArraySlice_l173_250_5);
  assign _zz_when_ArraySlice_l173_250_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_250_7);
  assign _zz_when_ArraySlice_l173_250_5 = {1'd0, _zz_when_ArraySlice_l173_250_6};
  assign _zz_when_ArraySlice_l173_250_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_250_7 = {1'd0, _zz_when_ArraySlice_l173_250_8};
  assign _zz_when_ArraySlice_l173_250_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_251 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_251_1);
  assign _zz_when_ArraySlice_l165_251_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_251_1 = {1'd0, _zz_when_ArraySlice_l165_251_2};
  assign _zz_when_ArraySlice_l166_251 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_251_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_251_2);
  assign _zz_when_ArraySlice_l166_251_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_251_3);
  assign _zz_when_ArraySlice_l166_251_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_251_3 = {1'd0, _zz_when_ArraySlice_l166_251_4};
  assign _zz__zz_when_ArraySlice_l112_251 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_251 = (_zz_when_ArraySlice_l113_251_1 - _zz_when_ArraySlice_l113_251_4);
  assign _zz_when_ArraySlice_l113_251_1 = (_zz_when_ArraySlice_l113_251_2 + _zz_when_ArraySlice_l113_251_3);
  assign _zz_when_ArraySlice_l113_251_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_251_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_251_4 = {1'd0, _zz_when_ArraySlice_l112_251};
  assign _zz__zz_when_ArraySlice_l173_251 = (_zz__zz_when_ArraySlice_l173_251_1 + _zz__zz_when_ArraySlice_l173_251_2);
  assign _zz__zz_when_ArraySlice_l173_251_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_251_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_251_3 = {1'd0, _zz_when_ArraySlice_l112_251};
  assign _zz_when_ArraySlice_l118_251_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_251 = _zz_when_ArraySlice_l118_251_1[5:0];
  assign _zz_when_ArraySlice_l173_251_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_251_1 = {1'd0, _zz_when_ArraySlice_l173_251_2};
  assign _zz_when_ArraySlice_l173_251_3 = (_zz_when_ArraySlice_l173_251_4 + _zz_when_ArraySlice_l173_251_9);
  assign _zz_when_ArraySlice_l173_251_4 = (_zz_when_ArraySlice_l173_251 - _zz_when_ArraySlice_l173_251_5);
  assign _zz_when_ArraySlice_l173_251_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_251_7);
  assign _zz_when_ArraySlice_l173_251_5 = {1'd0, _zz_when_ArraySlice_l173_251_6};
  assign _zz_when_ArraySlice_l173_251_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_251_7 = {1'd0, _zz_when_ArraySlice_l173_251_8};
  assign _zz_when_ArraySlice_l173_251_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_252 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_252_1);
  assign _zz_when_ArraySlice_l165_252_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_252 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_252_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_252_2);
  assign _zz_when_ArraySlice_l166_252_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_252_3);
  assign _zz_when_ArraySlice_l166_252_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_252 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_252 = (_zz_when_ArraySlice_l113_252_1 - _zz_when_ArraySlice_l113_252_4);
  assign _zz_when_ArraySlice_l113_252_1 = (_zz_when_ArraySlice_l113_252_2 + _zz_when_ArraySlice_l113_252_3);
  assign _zz_when_ArraySlice_l113_252_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_252_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_252_4 = {1'd0, _zz_when_ArraySlice_l112_252};
  assign _zz__zz_when_ArraySlice_l173_252 = (_zz__zz_when_ArraySlice_l173_252_1 + _zz__zz_when_ArraySlice_l173_252_2);
  assign _zz__zz_when_ArraySlice_l173_252_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_252_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_252_3 = {1'd0, _zz_when_ArraySlice_l112_252};
  assign _zz_when_ArraySlice_l118_252_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_252 = _zz_when_ArraySlice_l118_252_1[5:0];
  assign _zz_when_ArraySlice_l173_252_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_252_1 = {1'd0, _zz_when_ArraySlice_l173_252_2};
  assign _zz_when_ArraySlice_l173_252_3 = (_zz_when_ArraySlice_l173_252_4 + _zz_when_ArraySlice_l173_252_8);
  assign _zz_when_ArraySlice_l173_252_4 = (_zz_when_ArraySlice_l173_252 - _zz_when_ArraySlice_l173_252_5);
  assign _zz_when_ArraySlice_l173_252_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_252_7);
  assign _zz_when_ArraySlice_l173_252_5 = {1'd0, _zz_when_ArraySlice_l173_252_6};
  assign _zz_when_ArraySlice_l173_252_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_252_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_253 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_253_1);
  assign _zz_when_ArraySlice_l165_253_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_253_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_253 = {1'd0, _zz_when_ArraySlice_l166_253_1};
  assign _zz_when_ArraySlice_l166_253_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_253_3);
  assign _zz_when_ArraySlice_l166_253_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_253_4);
  assign _zz_when_ArraySlice_l166_253_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_253 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_253 = (_zz_when_ArraySlice_l113_253_1 - _zz_when_ArraySlice_l113_253_4);
  assign _zz_when_ArraySlice_l113_253_1 = (_zz_when_ArraySlice_l113_253_2 + _zz_when_ArraySlice_l113_253_3);
  assign _zz_when_ArraySlice_l113_253_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_253_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_253_4 = {1'd0, _zz_when_ArraySlice_l112_253};
  assign _zz__zz_when_ArraySlice_l173_253 = (_zz__zz_when_ArraySlice_l173_253_1 + _zz__zz_when_ArraySlice_l173_253_2);
  assign _zz__zz_when_ArraySlice_l173_253_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_253_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_253_3 = {1'd0, _zz_when_ArraySlice_l112_253};
  assign _zz_when_ArraySlice_l118_253_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_253 = _zz_when_ArraySlice_l118_253_1[5:0];
  assign _zz_when_ArraySlice_l173_253_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_253_1 = {2'd0, _zz_when_ArraySlice_l173_253_2};
  assign _zz_when_ArraySlice_l173_253_3 = (_zz_when_ArraySlice_l173_253_4 + _zz_when_ArraySlice_l173_253_8);
  assign _zz_when_ArraySlice_l173_253_4 = (_zz_when_ArraySlice_l173_253 - _zz_when_ArraySlice_l173_253_5);
  assign _zz_when_ArraySlice_l173_253_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_253_7);
  assign _zz_when_ArraySlice_l173_253_5 = {1'd0, _zz_when_ArraySlice_l173_253_6};
  assign _zz_when_ArraySlice_l173_253_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_253_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_254 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_254_1);
  assign _zz_when_ArraySlice_l165_254_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_254_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_254 = {1'd0, _zz_when_ArraySlice_l166_254_1};
  assign _zz_when_ArraySlice_l166_254_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_254_3);
  assign _zz_when_ArraySlice_l166_254_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_254_4);
  assign _zz_when_ArraySlice_l166_254_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_254 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_254 = (_zz_when_ArraySlice_l113_254_1 - _zz_when_ArraySlice_l113_254_4);
  assign _zz_when_ArraySlice_l113_254_1 = (_zz_when_ArraySlice_l113_254_2 + _zz_when_ArraySlice_l113_254_3);
  assign _zz_when_ArraySlice_l113_254_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_254_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_254_4 = {1'd0, _zz_when_ArraySlice_l112_254};
  assign _zz__zz_when_ArraySlice_l173_254 = (_zz__zz_when_ArraySlice_l173_254_1 + _zz__zz_when_ArraySlice_l173_254_2);
  assign _zz__zz_when_ArraySlice_l173_254_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_254_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_254_3 = {1'd0, _zz_when_ArraySlice_l112_254};
  assign _zz_when_ArraySlice_l118_254_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_254 = _zz_when_ArraySlice_l118_254_1[5:0];
  assign _zz_when_ArraySlice_l173_254_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_254_1 = {2'd0, _zz_when_ArraySlice_l173_254_2};
  assign _zz_when_ArraySlice_l173_254_3 = (_zz_when_ArraySlice_l173_254_4 + _zz_when_ArraySlice_l173_254_8);
  assign _zz_when_ArraySlice_l173_254_4 = (_zz_when_ArraySlice_l173_254 - _zz_when_ArraySlice_l173_254_5);
  assign _zz_when_ArraySlice_l173_254_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_254_7);
  assign _zz_when_ArraySlice_l173_254_5 = {1'd0, _zz_when_ArraySlice_l173_254_6};
  assign _zz_when_ArraySlice_l173_254_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_254_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_255 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_255_1);
  assign _zz_when_ArraySlice_l165_255_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_255_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_255 = {2'd0, _zz_when_ArraySlice_l166_255_1};
  assign _zz_when_ArraySlice_l166_255_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_255_3);
  assign _zz_when_ArraySlice_l166_255_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_255_4);
  assign _zz_when_ArraySlice_l166_255_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_255 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_255 = (_zz_when_ArraySlice_l113_255_1 - _zz_when_ArraySlice_l113_255_4);
  assign _zz_when_ArraySlice_l113_255_1 = (_zz_when_ArraySlice_l113_255_2 + _zz_when_ArraySlice_l113_255_3);
  assign _zz_when_ArraySlice_l113_255_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_255_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_255_4 = {1'd0, _zz_when_ArraySlice_l112_255};
  assign _zz__zz_when_ArraySlice_l173_255 = (_zz__zz_when_ArraySlice_l173_255_1 + _zz__zz_when_ArraySlice_l173_255_2);
  assign _zz__zz_when_ArraySlice_l173_255_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_255_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_255_3 = {1'd0, _zz_when_ArraySlice_l112_255};
  assign _zz_when_ArraySlice_l118_255_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_255 = _zz_when_ArraySlice_l118_255_1[5:0];
  assign _zz_when_ArraySlice_l173_255_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_255_1 = {3'd0, _zz_when_ArraySlice_l173_255_2};
  assign _zz_when_ArraySlice_l173_255_3 = (_zz_when_ArraySlice_l173_255_4 + _zz_when_ArraySlice_l173_255_8);
  assign _zz_when_ArraySlice_l173_255_4 = (_zz_when_ArraySlice_l173_255 - _zz_when_ArraySlice_l173_255_5);
  assign _zz_when_ArraySlice_l173_255_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_255_7);
  assign _zz_when_ArraySlice_l173_255_5 = {1'd0, _zz_when_ArraySlice_l173_255_6};
  assign _zz_when_ArraySlice_l173_255_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_255_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_1_63 = 1'b1;
  assign _zz_selectReadFifo_1_62 = {5'd0, _zz_selectReadFifo_1_63};
  assign _zz_when_ArraySlice_l315_1_1 = (_zz_when_ArraySlice_l315_1_2 % aReg);
  assign _zz_when_ArraySlice_l315_1_2 = (handshakeTimes_1_value + _zz_when_ArraySlice_l315_1_3);
  assign _zz_when_ArraySlice_l315_1_4 = 1'b1;
  assign _zz_when_ArraySlice_l315_1_3 = {12'd0, _zz_when_ArraySlice_l315_1_4};
  assign _zz_when_ArraySlice_l301_1_1 = (selectReadFifo_1 + _zz_when_ArraySlice_l301_1_2);
  assign _zz_when_ArraySlice_l301_1_3 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l301_1_2 = {2'd0, _zz_when_ArraySlice_l301_1_3};
  assign _zz_when_ArraySlice_l322_1_2 = (_zz_when_ArraySlice_l322_1_3 - _zz_when_ArraySlice_l322_1_4);
  assign _zz_when_ArraySlice_l322_1_1 = {7'd0, _zz_when_ArraySlice_l322_1_2};
  assign _zz_when_ArraySlice_l322_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l322_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l322_1_4 = {5'd0, _zz_when_ArraySlice_l322_1_5};
  assign _zz_when_ArraySlice_l240_2_1 = (selectReadFifo_2 + _zz_when_ArraySlice_l240_2_2);
  assign _zz_when_ArraySlice_l240_2_3 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l240_2_2 = {1'd0, _zz_when_ArraySlice_l240_2_3};
  assign _zz_when_ArraySlice_l241_2_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l241_2_3);
  assign _zz_when_ArraySlice_l241_2_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l241_2_3 = {1'd0, _zz_when_ArraySlice_l241_2_4};
  assign _zz__zz_outputStreamArrayData_2_valid_1_2 = (bReg * 2'b10);
  assign _zz__zz_outputStreamArrayData_2_valid_1_1 = {1'd0, _zz__zz_outputStreamArrayData_2_valid_1_2};
  assign _zz_when_ArraySlice_l247_2_2 = 1'b1;
  assign _zz_when_ArraySlice_l247_2_1 = {6'd0, _zz_when_ArraySlice_l247_2_2};
  assign _zz_when_ArraySlice_l247_2_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l247_2_5);
  assign _zz_when_ArraySlice_l247_2_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l247_2_5 = {1'd0, _zz_when_ArraySlice_l247_2_6};
  assign _zz_when_ArraySlice_l248_2_2 = (_zz_when_ArraySlice_l248_2_3 - _zz_when_ArraySlice_l248_2_4);
  assign _zz_when_ArraySlice_l248_2_1 = {7'd0, _zz_when_ArraySlice_l248_2_2};
  assign _zz_when_ArraySlice_l248_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l248_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l248_2_4 = {5'd0, _zz_when_ArraySlice_l248_2_5};
  assign _zz_selectReadFifo_2_32 = (selectReadFifo_2 - _zz_selectReadFifo_2_33);
  assign _zz_selectReadFifo_2_33 = {3'd0, bReg};
  assign _zz_selectReadFifo_2_35 = 1'b1;
  assign _zz_selectReadFifo_2_34 = {5'd0, _zz_selectReadFifo_2_35};
  assign _zz_selectReadFifo_2_37 = 1'b1;
  assign _zz_selectReadFifo_2_36 = {5'd0, _zz_selectReadFifo_2_37};
  assign _zz_when_ArraySlice_l251_2_1 = (_zz_when_ArraySlice_l251_2_2 % aReg);
  assign _zz_when_ArraySlice_l251_2_2 = (handshakeTimes_2_value + _zz_when_ArraySlice_l251_2_3);
  assign _zz_when_ArraySlice_l251_2_4 = 1'b1;
  assign _zz_when_ArraySlice_l251_2_3 = {12'd0, _zz_when_ArraySlice_l251_2_4};
  assign _zz_when_ArraySlice_l256_2_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l256_2_3);
  assign _zz_when_ArraySlice_l256_2_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l256_2_3 = {1'd0, _zz_when_ArraySlice_l256_2_4};
  assign _zz_when_ArraySlice_l256_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l256_2_5 = {6'd0, _zz_when_ArraySlice_l256_2_6};
  assign _zz_when_ArraySlice_l257_2_2 = (_zz_when_ArraySlice_l257_2_3 - _zz_when_ArraySlice_l257_2_4);
  assign _zz_when_ArraySlice_l257_2_1 = {7'd0, _zz_when_ArraySlice_l257_2_2};
  assign _zz_when_ArraySlice_l257_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l257_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l257_2_4 = {5'd0, _zz_when_ArraySlice_l257_2_5};
  assign _zz__zz_when_ArraySlice_l94_30 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_30 = (_zz_when_ArraySlice_l95_30_1 - _zz_when_ArraySlice_l95_30_4);
  assign _zz_when_ArraySlice_l95_30_1 = (_zz_when_ArraySlice_l95_30_2 + _zz_when_ArraySlice_l95_30_3);
  assign _zz_when_ArraySlice_l95_30_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_30_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_30_4 = {1'd0, _zz_when_ArraySlice_l94_30};
  assign _zz__zz_when_ArraySlice_l259_2_1 = (_zz__zz_when_ArraySlice_l259_2_2 + _zz__zz_when_ArraySlice_l259_2_3);
  assign _zz__zz_when_ArraySlice_l259_2_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l259_2_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l259_2_4 = {1'd0, _zz_when_ArraySlice_l94_30};
  assign _zz_when_ArraySlice_l99_30_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_30 = _zz_when_ArraySlice_l99_30_1[5:0];
  assign _zz_when_ArraySlice_l259_2_1 = (outSliceNumb_2_value + _zz_when_ArraySlice_l259_2_2);
  assign _zz_when_ArraySlice_l259_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l259_2_2 = {6'd0, _zz_when_ArraySlice_l259_2_3};
  assign _zz_when_ArraySlice_l259_2_4 = (_zz_when_ArraySlice_l259_2 / aReg);
  assign _zz_selectReadFifo_2_38 = (selectReadFifo_2 - _zz_selectReadFifo_2_39);
  assign _zz_selectReadFifo_2_39 = {3'd0, bReg};
  assign _zz_selectReadFifo_2_41 = 1'b1;
  assign _zz_selectReadFifo_2_40 = {5'd0, _zz_selectReadFifo_2_41};
  assign _zz_selectReadFifo_2_42 = (selectReadFifo_2 + _zz_selectReadFifo_2_43);
  assign _zz_selectReadFifo_2_43 = (3'b111 * bReg);
  assign _zz_selectReadFifo_2_45 = 1'b1;
  assign _zz_selectReadFifo_2_44 = {5'd0, _zz_selectReadFifo_2_45};
  assign _zz_when_ArraySlice_l165_256 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_256_1);
  assign _zz_when_ArraySlice_l165_256_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_256_1 = {3'd0, _zz_when_ArraySlice_l165_256_2};
  assign _zz_when_ArraySlice_l166_256 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_256_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_256_3);
  assign _zz_when_ArraySlice_l166_256_1 = {1'd0, _zz_when_ArraySlice_l166_256_2};
  assign _zz_when_ArraySlice_l166_256_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_256_4);
  assign _zz_when_ArraySlice_l166_256_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_256_4 = {3'd0, _zz_when_ArraySlice_l166_256_5};
  assign _zz__zz_when_ArraySlice_l112_256 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_256 = (_zz_when_ArraySlice_l113_256_1 - _zz_when_ArraySlice_l113_256_4);
  assign _zz_when_ArraySlice_l113_256_1 = (_zz_when_ArraySlice_l113_256_2 + _zz_when_ArraySlice_l113_256_3);
  assign _zz_when_ArraySlice_l113_256_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_256_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_256_4 = {1'd0, _zz_when_ArraySlice_l112_256};
  assign _zz__zz_when_ArraySlice_l173_256 = (_zz__zz_when_ArraySlice_l173_256_1 + _zz__zz_when_ArraySlice_l173_256_2);
  assign _zz__zz_when_ArraySlice_l173_256_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_256_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_256_3 = {1'd0, _zz_when_ArraySlice_l112_256};
  assign _zz_when_ArraySlice_l118_256_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_256 = _zz_when_ArraySlice_l118_256_1[5:0];
  assign _zz_when_ArraySlice_l173_256_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_256_2 = (_zz_when_ArraySlice_l173_256_3 + _zz_when_ArraySlice_l173_256_8);
  assign _zz_when_ArraySlice_l173_256_3 = (_zz_when_ArraySlice_l173_256 - _zz_when_ArraySlice_l173_256_4);
  assign _zz_when_ArraySlice_l173_256_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_256_6);
  assign _zz_when_ArraySlice_l173_256_4 = {1'd0, _zz_when_ArraySlice_l173_256_5};
  assign _zz_when_ArraySlice_l173_256_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_256_6 = {3'd0, _zz_when_ArraySlice_l173_256_7};
  assign _zz_when_ArraySlice_l173_256_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_257 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_257_1);
  assign _zz_when_ArraySlice_l165_257_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_257_1 = {2'd0, _zz_when_ArraySlice_l165_257_2};
  assign _zz_when_ArraySlice_l166_257 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_257_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_257_2);
  assign _zz_when_ArraySlice_l166_257_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_257_3);
  assign _zz_when_ArraySlice_l166_257_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_257_3 = {2'd0, _zz_when_ArraySlice_l166_257_4};
  assign _zz__zz_when_ArraySlice_l112_257 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_257 = (_zz_when_ArraySlice_l113_257_1 - _zz_when_ArraySlice_l113_257_4);
  assign _zz_when_ArraySlice_l113_257_1 = (_zz_when_ArraySlice_l113_257_2 + _zz_when_ArraySlice_l113_257_3);
  assign _zz_when_ArraySlice_l113_257_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_257_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_257_4 = {1'd0, _zz_when_ArraySlice_l112_257};
  assign _zz__zz_when_ArraySlice_l173_257 = (_zz__zz_when_ArraySlice_l173_257_1 + _zz__zz_when_ArraySlice_l173_257_2);
  assign _zz__zz_when_ArraySlice_l173_257_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_257_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_257_3 = {1'd0, _zz_when_ArraySlice_l112_257};
  assign _zz_when_ArraySlice_l118_257_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_257 = _zz_when_ArraySlice_l118_257_1[5:0];
  assign _zz_when_ArraySlice_l173_257_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_257_1 = {1'd0, _zz_when_ArraySlice_l173_257_2};
  assign _zz_when_ArraySlice_l173_257_3 = (_zz_when_ArraySlice_l173_257_4 + _zz_when_ArraySlice_l173_257_9);
  assign _zz_when_ArraySlice_l173_257_4 = (_zz_when_ArraySlice_l173_257 - _zz_when_ArraySlice_l173_257_5);
  assign _zz_when_ArraySlice_l173_257_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_257_7);
  assign _zz_when_ArraySlice_l173_257_5 = {1'd0, _zz_when_ArraySlice_l173_257_6};
  assign _zz_when_ArraySlice_l173_257_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_257_7 = {2'd0, _zz_when_ArraySlice_l173_257_8};
  assign _zz_when_ArraySlice_l173_257_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_258 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_258_1);
  assign _zz_when_ArraySlice_l165_258_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_258_1 = {1'd0, _zz_when_ArraySlice_l165_258_2};
  assign _zz_when_ArraySlice_l166_258 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_258_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_258_2);
  assign _zz_when_ArraySlice_l166_258_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_258_3);
  assign _zz_when_ArraySlice_l166_258_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_258_3 = {1'd0, _zz_when_ArraySlice_l166_258_4};
  assign _zz__zz_when_ArraySlice_l112_258 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_258 = (_zz_when_ArraySlice_l113_258_1 - _zz_when_ArraySlice_l113_258_4);
  assign _zz_when_ArraySlice_l113_258_1 = (_zz_when_ArraySlice_l113_258_2 + _zz_when_ArraySlice_l113_258_3);
  assign _zz_when_ArraySlice_l113_258_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_258_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_258_4 = {1'd0, _zz_when_ArraySlice_l112_258};
  assign _zz__zz_when_ArraySlice_l173_258 = (_zz__zz_when_ArraySlice_l173_258_1 + _zz__zz_when_ArraySlice_l173_258_2);
  assign _zz__zz_when_ArraySlice_l173_258_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_258_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_258_3 = {1'd0, _zz_when_ArraySlice_l112_258};
  assign _zz_when_ArraySlice_l118_258_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_258 = _zz_when_ArraySlice_l118_258_1[5:0];
  assign _zz_when_ArraySlice_l173_258_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_258_1 = {1'd0, _zz_when_ArraySlice_l173_258_2};
  assign _zz_when_ArraySlice_l173_258_3 = (_zz_when_ArraySlice_l173_258_4 + _zz_when_ArraySlice_l173_258_9);
  assign _zz_when_ArraySlice_l173_258_4 = (_zz_when_ArraySlice_l173_258 - _zz_when_ArraySlice_l173_258_5);
  assign _zz_when_ArraySlice_l173_258_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_258_7);
  assign _zz_when_ArraySlice_l173_258_5 = {1'd0, _zz_when_ArraySlice_l173_258_6};
  assign _zz_when_ArraySlice_l173_258_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_258_7 = {1'd0, _zz_when_ArraySlice_l173_258_8};
  assign _zz_when_ArraySlice_l173_258_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_259 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_259_1);
  assign _zz_when_ArraySlice_l165_259_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_259_1 = {1'd0, _zz_when_ArraySlice_l165_259_2};
  assign _zz_when_ArraySlice_l166_259 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_259_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_259_2);
  assign _zz_when_ArraySlice_l166_259_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_259_3);
  assign _zz_when_ArraySlice_l166_259_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_259_3 = {1'd0, _zz_when_ArraySlice_l166_259_4};
  assign _zz__zz_when_ArraySlice_l112_259 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_259 = (_zz_when_ArraySlice_l113_259_1 - _zz_when_ArraySlice_l113_259_4);
  assign _zz_when_ArraySlice_l113_259_1 = (_zz_when_ArraySlice_l113_259_2 + _zz_when_ArraySlice_l113_259_3);
  assign _zz_when_ArraySlice_l113_259_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_259_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_259_4 = {1'd0, _zz_when_ArraySlice_l112_259};
  assign _zz__zz_when_ArraySlice_l173_259 = (_zz__zz_when_ArraySlice_l173_259_1 + _zz__zz_when_ArraySlice_l173_259_2);
  assign _zz__zz_when_ArraySlice_l173_259_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_259_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_259_3 = {1'd0, _zz_when_ArraySlice_l112_259};
  assign _zz_when_ArraySlice_l118_259_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_259 = _zz_when_ArraySlice_l118_259_1[5:0];
  assign _zz_when_ArraySlice_l173_259_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_259_1 = {1'd0, _zz_when_ArraySlice_l173_259_2};
  assign _zz_when_ArraySlice_l173_259_3 = (_zz_when_ArraySlice_l173_259_4 + _zz_when_ArraySlice_l173_259_9);
  assign _zz_when_ArraySlice_l173_259_4 = (_zz_when_ArraySlice_l173_259 - _zz_when_ArraySlice_l173_259_5);
  assign _zz_when_ArraySlice_l173_259_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_259_7);
  assign _zz_when_ArraySlice_l173_259_5 = {1'd0, _zz_when_ArraySlice_l173_259_6};
  assign _zz_when_ArraySlice_l173_259_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_259_7 = {1'd0, _zz_when_ArraySlice_l173_259_8};
  assign _zz_when_ArraySlice_l173_259_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_260 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_260_1);
  assign _zz_when_ArraySlice_l165_260_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_260 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_260_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_260_2);
  assign _zz_when_ArraySlice_l166_260_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_260_3);
  assign _zz_when_ArraySlice_l166_260_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_260 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_260 = (_zz_when_ArraySlice_l113_260_1 - _zz_when_ArraySlice_l113_260_4);
  assign _zz_when_ArraySlice_l113_260_1 = (_zz_when_ArraySlice_l113_260_2 + _zz_when_ArraySlice_l113_260_3);
  assign _zz_when_ArraySlice_l113_260_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_260_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_260_4 = {1'd0, _zz_when_ArraySlice_l112_260};
  assign _zz__zz_when_ArraySlice_l173_260 = (_zz__zz_when_ArraySlice_l173_260_1 + _zz__zz_when_ArraySlice_l173_260_2);
  assign _zz__zz_when_ArraySlice_l173_260_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_260_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_260_3 = {1'd0, _zz_when_ArraySlice_l112_260};
  assign _zz_when_ArraySlice_l118_260_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_260 = _zz_when_ArraySlice_l118_260_1[5:0];
  assign _zz_when_ArraySlice_l173_260_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_260_1 = {1'd0, _zz_when_ArraySlice_l173_260_2};
  assign _zz_when_ArraySlice_l173_260_3 = (_zz_when_ArraySlice_l173_260_4 + _zz_when_ArraySlice_l173_260_8);
  assign _zz_when_ArraySlice_l173_260_4 = (_zz_when_ArraySlice_l173_260 - _zz_when_ArraySlice_l173_260_5);
  assign _zz_when_ArraySlice_l173_260_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_260_7);
  assign _zz_when_ArraySlice_l173_260_5 = {1'd0, _zz_when_ArraySlice_l173_260_6};
  assign _zz_when_ArraySlice_l173_260_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_260_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_261 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_261_1);
  assign _zz_when_ArraySlice_l165_261_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_261_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_261 = {1'd0, _zz_when_ArraySlice_l166_261_1};
  assign _zz_when_ArraySlice_l166_261_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_261_3);
  assign _zz_when_ArraySlice_l166_261_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_261_4);
  assign _zz_when_ArraySlice_l166_261_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_261 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_261 = (_zz_when_ArraySlice_l113_261_1 - _zz_when_ArraySlice_l113_261_4);
  assign _zz_when_ArraySlice_l113_261_1 = (_zz_when_ArraySlice_l113_261_2 + _zz_when_ArraySlice_l113_261_3);
  assign _zz_when_ArraySlice_l113_261_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_261_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_261_4 = {1'd0, _zz_when_ArraySlice_l112_261};
  assign _zz__zz_when_ArraySlice_l173_261 = (_zz__zz_when_ArraySlice_l173_261_1 + _zz__zz_when_ArraySlice_l173_261_2);
  assign _zz__zz_when_ArraySlice_l173_261_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_261_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_261_3 = {1'd0, _zz_when_ArraySlice_l112_261};
  assign _zz_when_ArraySlice_l118_261_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_261 = _zz_when_ArraySlice_l118_261_1[5:0];
  assign _zz_when_ArraySlice_l173_261_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_261_1 = {2'd0, _zz_when_ArraySlice_l173_261_2};
  assign _zz_when_ArraySlice_l173_261_3 = (_zz_when_ArraySlice_l173_261_4 + _zz_when_ArraySlice_l173_261_8);
  assign _zz_when_ArraySlice_l173_261_4 = (_zz_when_ArraySlice_l173_261 - _zz_when_ArraySlice_l173_261_5);
  assign _zz_when_ArraySlice_l173_261_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_261_7);
  assign _zz_when_ArraySlice_l173_261_5 = {1'd0, _zz_when_ArraySlice_l173_261_6};
  assign _zz_when_ArraySlice_l173_261_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_261_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_262 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_262_1);
  assign _zz_when_ArraySlice_l165_262_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_262_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_262 = {1'd0, _zz_when_ArraySlice_l166_262_1};
  assign _zz_when_ArraySlice_l166_262_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_262_3);
  assign _zz_when_ArraySlice_l166_262_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_262_4);
  assign _zz_when_ArraySlice_l166_262_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_262 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_262 = (_zz_when_ArraySlice_l113_262_1 - _zz_when_ArraySlice_l113_262_4);
  assign _zz_when_ArraySlice_l113_262_1 = (_zz_when_ArraySlice_l113_262_2 + _zz_when_ArraySlice_l113_262_3);
  assign _zz_when_ArraySlice_l113_262_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_262_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_262_4 = {1'd0, _zz_when_ArraySlice_l112_262};
  assign _zz__zz_when_ArraySlice_l173_262 = (_zz__zz_when_ArraySlice_l173_262_1 + _zz__zz_when_ArraySlice_l173_262_2);
  assign _zz__zz_when_ArraySlice_l173_262_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_262_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_262_3 = {1'd0, _zz_when_ArraySlice_l112_262};
  assign _zz_when_ArraySlice_l118_262_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_262 = _zz_when_ArraySlice_l118_262_1[5:0];
  assign _zz_when_ArraySlice_l173_262_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_262_1 = {2'd0, _zz_when_ArraySlice_l173_262_2};
  assign _zz_when_ArraySlice_l173_262_3 = (_zz_when_ArraySlice_l173_262_4 + _zz_when_ArraySlice_l173_262_8);
  assign _zz_when_ArraySlice_l173_262_4 = (_zz_when_ArraySlice_l173_262 - _zz_when_ArraySlice_l173_262_5);
  assign _zz_when_ArraySlice_l173_262_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_262_7);
  assign _zz_when_ArraySlice_l173_262_5 = {1'd0, _zz_when_ArraySlice_l173_262_6};
  assign _zz_when_ArraySlice_l173_262_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_262_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_263 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_263_1);
  assign _zz_when_ArraySlice_l165_263_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_263_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_263 = {2'd0, _zz_when_ArraySlice_l166_263_1};
  assign _zz_when_ArraySlice_l166_263_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_263_3);
  assign _zz_when_ArraySlice_l166_263_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_263_4);
  assign _zz_when_ArraySlice_l166_263_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_263 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_263 = (_zz_when_ArraySlice_l113_263_1 - _zz_when_ArraySlice_l113_263_4);
  assign _zz_when_ArraySlice_l113_263_1 = (_zz_when_ArraySlice_l113_263_2 + _zz_when_ArraySlice_l113_263_3);
  assign _zz_when_ArraySlice_l113_263_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_263_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_263_4 = {1'd0, _zz_when_ArraySlice_l112_263};
  assign _zz__zz_when_ArraySlice_l173_263 = (_zz__zz_when_ArraySlice_l173_263_1 + _zz__zz_when_ArraySlice_l173_263_2);
  assign _zz__zz_when_ArraySlice_l173_263_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_263_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_263_3 = {1'd0, _zz_when_ArraySlice_l112_263};
  assign _zz_when_ArraySlice_l118_263_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_263 = _zz_when_ArraySlice_l118_263_1[5:0];
  assign _zz_when_ArraySlice_l173_263_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_263_1 = {3'd0, _zz_when_ArraySlice_l173_263_2};
  assign _zz_when_ArraySlice_l173_263_3 = (_zz_when_ArraySlice_l173_263_4 + _zz_when_ArraySlice_l173_263_8);
  assign _zz_when_ArraySlice_l173_263_4 = (_zz_when_ArraySlice_l173_263 - _zz_when_ArraySlice_l173_263_5);
  assign _zz_when_ArraySlice_l173_263_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_263_7);
  assign _zz_when_ArraySlice_l173_263_5 = {1'd0, _zz_when_ArraySlice_l173_263_6};
  assign _zz_when_ArraySlice_l173_263_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_263_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l268_2_1 = (_zz_when_ArraySlice_l268_2_2 + _zz_when_ArraySlice_l268_2_7);
  assign _zz_when_ArraySlice_l268_2_2 = (_zz_when_ArraySlice_l268_2_3 + _zz_when_ArraySlice_l268_2_5);
  assign _zz_when_ArraySlice_l268_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l268_2_4);
  assign _zz_when_ArraySlice_l268_2_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l268_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l268_2_5 = {5'd0, _zz_when_ArraySlice_l268_2_6};
  assign _zz_when_ArraySlice_l268_2_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l268_2_7 = {1'd0, _zz_when_ArraySlice_l268_2_8};
  assign _zz_selectReadFifo_2_47 = 1'b1;
  assign _zz_selectReadFifo_2_46 = {5'd0, _zz_selectReadFifo_2_47};
  assign _zz_when_ArraySlice_l272_2_1 = (_zz_when_ArraySlice_l272_2_2 % aReg);
  assign _zz_when_ArraySlice_l272_2_2 = (handshakeTimes_2_value + _zz_when_ArraySlice_l272_2_3);
  assign _zz_when_ArraySlice_l272_2_4 = 1'b1;
  assign _zz_when_ArraySlice_l272_2_3 = {12'd0, _zz_when_ArraySlice_l272_2_4};
  assign _zz_when_ArraySlice_l276_2_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l276_2_3);
  assign _zz_when_ArraySlice_l276_2_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l276_2_3 = {1'd0, _zz_when_ArraySlice_l276_2_4};
  assign _zz_when_ArraySlice_l277_2_2 = (_zz_when_ArraySlice_l277_2_3 - _zz_when_ArraySlice_l277_2_4);
  assign _zz_when_ArraySlice_l277_2_1 = {7'd0, _zz_when_ArraySlice_l277_2_2};
  assign _zz_when_ArraySlice_l277_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l277_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l277_2_4 = {5'd0, _zz_when_ArraySlice_l277_2_5};
  assign _zz__zz_when_ArraySlice_l94_31 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_31 = (_zz_when_ArraySlice_l95_31_1 - _zz_when_ArraySlice_l95_31_4);
  assign _zz_when_ArraySlice_l95_31_1 = (_zz_when_ArraySlice_l95_31_2 + _zz_when_ArraySlice_l95_31_3);
  assign _zz_when_ArraySlice_l95_31_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_31_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_31_4 = {1'd0, _zz_when_ArraySlice_l94_31};
  assign _zz__zz_when_ArraySlice_l279_2_1 = (_zz__zz_when_ArraySlice_l279_2_2 + _zz__zz_when_ArraySlice_l279_2_3);
  assign _zz__zz_when_ArraySlice_l279_2_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l279_2_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l279_2_4 = {1'd0, _zz_when_ArraySlice_l94_31};
  assign _zz_when_ArraySlice_l99_31_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_31 = _zz_when_ArraySlice_l99_31_1[5:0];
  assign _zz_when_ArraySlice_l279_2_1 = (outSliceNumb_2_value + _zz_when_ArraySlice_l279_2_2);
  assign _zz_when_ArraySlice_l279_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l279_2_2 = {6'd0, _zz_when_ArraySlice_l279_2_3};
  assign _zz_when_ArraySlice_l279_2_4 = (_zz_when_ArraySlice_l279_2 / aReg);
  assign _zz_selectReadFifo_2_48 = (selectReadFifo_2 - _zz_selectReadFifo_2_49);
  assign _zz_selectReadFifo_2_49 = {3'd0, bReg};
  assign _zz_selectReadFifo_2_51 = 1'b1;
  assign _zz_selectReadFifo_2_50 = {5'd0, _zz_selectReadFifo_2_51};
  assign _zz_selectReadFifo_2_52 = (selectReadFifo_2 + _zz_selectReadFifo_2_53);
  assign _zz_selectReadFifo_2_53 = (3'b111 * bReg);
  assign _zz_selectReadFifo_2_55 = 1'b1;
  assign _zz_selectReadFifo_2_54 = {5'd0, _zz_selectReadFifo_2_55};
  assign _zz_when_ArraySlice_l165_264 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_264_1);
  assign _zz_when_ArraySlice_l165_264_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_264_1 = {3'd0, _zz_when_ArraySlice_l165_264_2};
  assign _zz_when_ArraySlice_l166_264 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_264_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_264_3);
  assign _zz_when_ArraySlice_l166_264_1 = {1'd0, _zz_when_ArraySlice_l166_264_2};
  assign _zz_when_ArraySlice_l166_264_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_264_4);
  assign _zz_when_ArraySlice_l166_264_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_264_4 = {3'd0, _zz_when_ArraySlice_l166_264_5};
  assign _zz__zz_when_ArraySlice_l112_264 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_264 = (_zz_when_ArraySlice_l113_264_1 - _zz_when_ArraySlice_l113_264_4);
  assign _zz_when_ArraySlice_l113_264_1 = (_zz_when_ArraySlice_l113_264_2 + _zz_when_ArraySlice_l113_264_3);
  assign _zz_when_ArraySlice_l113_264_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_264_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_264_4 = {1'd0, _zz_when_ArraySlice_l112_264};
  assign _zz__zz_when_ArraySlice_l173_264 = (_zz__zz_when_ArraySlice_l173_264_1 + _zz__zz_when_ArraySlice_l173_264_2);
  assign _zz__zz_when_ArraySlice_l173_264_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_264_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_264_3 = {1'd0, _zz_when_ArraySlice_l112_264};
  assign _zz_when_ArraySlice_l118_264_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_264 = _zz_when_ArraySlice_l118_264_1[5:0];
  assign _zz_when_ArraySlice_l173_264_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_264_2 = (_zz_when_ArraySlice_l173_264_3 + _zz_when_ArraySlice_l173_264_8);
  assign _zz_when_ArraySlice_l173_264_3 = (_zz_when_ArraySlice_l173_264 - _zz_when_ArraySlice_l173_264_4);
  assign _zz_when_ArraySlice_l173_264_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_264_6);
  assign _zz_when_ArraySlice_l173_264_4 = {1'd0, _zz_when_ArraySlice_l173_264_5};
  assign _zz_when_ArraySlice_l173_264_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_264_6 = {3'd0, _zz_when_ArraySlice_l173_264_7};
  assign _zz_when_ArraySlice_l173_264_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_265 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_265_1);
  assign _zz_when_ArraySlice_l165_265_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_265_1 = {2'd0, _zz_when_ArraySlice_l165_265_2};
  assign _zz_when_ArraySlice_l166_265 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_265_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_265_2);
  assign _zz_when_ArraySlice_l166_265_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_265_3);
  assign _zz_when_ArraySlice_l166_265_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_265_3 = {2'd0, _zz_when_ArraySlice_l166_265_4};
  assign _zz__zz_when_ArraySlice_l112_265 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_265 = (_zz_when_ArraySlice_l113_265_1 - _zz_when_ArraySlice_l113_265_4);
  assign _zz_when_ArraySlice_l113_265_1 = (_zz_when_ArraySlice_l113_265_2 + _zz_when_ArraySlice_l113_265_3);
  assign _zz_when_ArraySlice_l113_265_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_265_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_265_4 = {1'd0, _zz_when_ArraySlice_l112_265};
  assign _zz__zz_when_ArraySlice_l173_265 = (_zz__zz_when_ArraySlice_l173_265_1 + _zz__zz_when_ArraySlice_l173_265_2);
  assign _zz__zz_when_ArraySlice_l173_265_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_265_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_265_3 = {1'd0, _zz_when_ArraySlice_l112_265};
  assign _zz_when_ArraySlice_l118_265_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_265 = _zz_when_ArraySlice_l118_265_1[5:0];
  assign _zz_when_ArraySlice_l173_265_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_265_1 = {1'd0, _zz_when_ArraySlice_l173_265_2};
  assign _zz_when_ArraySlice_l173_265_3 = (_zz_when_ArraySlice_l173_265_4 + _zz_when_ArraySlice_l173_265_9);
  assign _zz_when_ArraySlice_l173_265_4 = (_zz_when_ArraySlice_l173_265 - _zz_when_ArraySlice_l173_265_5);
  assign _zz_when_ArraySlice_l173_265_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_265_7);
  assign _zz_when_ArraySlice_l173_265_5 = {1'd0, _zz_when_ArraySlice_l173_265_6};
  assign _zz_when_ArraySlice_l173_265_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_265_7 = {2'd0, _zz_when_ArraySlice_l173_265_8};
  assign _zz_when_ArraySlice_l173_265_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_266 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_266_1);
  assign _zz_when_ArraySlice_l165_266_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_266_1 = {1'd0, _zz_when_ArraySlice_l165_266_2};
  assign _zz_when_ArraySlice_l166_266 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_266_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_266_2);
  assign _zz_when_ArraySlice_l166_266_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_266_3);
  assign _zz_when_ArraySlice_l166_266_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_266_3 = {1'd0, _zz_when_ArraySlice_l166_266_4};
  assign _zz__zz_when_ArraySlice_l112_266 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_266 = (_zz_when_ArraySlice_l113_266_1 - _zz_when_ArraySlice_l113_266_4);
  assign _zz_when_ArraySlice_l113_266_1 = (_zz_when_ArraySlice_l113_266_2 + _zz_when_ArraySlice_l113_266_3);
  assign _zz_when_ArraySlice_l113_266_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_266_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_266_4 = {1'd0, _zz_when_ArraySlice_l112_266};
  assign _zz__zz_when_ArraySlice_l173_266 = (_zz__zz_when_ArraySlice_l173_266_1 + _zz__zz_when_ArraySlice_l173_266_2);
  assign _zz__zz_when_ArraySlice_l173_266_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_266_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_266_3 = {1'd0, _zz_when_ArraySlice_l112_266};
  assign _zz_when_ArraySlice_l118_266_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_266 = _zz_when_ArraySlice_l118_266_1[5:0];
  assign _zz_when_ArraySlice_l173_266_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_266_1 = {1'd0, _zz_when_ArraySlice_l173_266_2};
  assign _zz_when_ArraySlice_l173_266_3 = (_zz_when_ArraySlice_l173_266_4 + _zz_when_ArraySlice_l173_266_9);
  assign _zz_when_ArraySlice_l173_266_4 = (_zz_when_ArraySlice_l173_266 - _zz_when_ArraySlice_l173_266_5);
  assign _zz_when_ArraySlice_l173_266_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_266_7);
  assign _zz_when_ArraySlice_l173_266_5 = {1'd0, _zz_when_ArraySlice_l173_266_6};
  assign _zz_when_ArraySlice_l173_266_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_266_7 = {1'd0, _zz_when_ArraySlice_l173_266_8};
  assign _zz_when_ArraySlice_l173_266_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_267 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_267_1);
  assign _zz_when_ArraySlice_l165_267_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_267_1 = {1'd0, _zz_when_ArraySlice_l165_267_2};
  assign _zz_when_ArraySlice_l166_267 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_267_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_267_2);
  assign _zz_when_ArraySlice_l166_267_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_267_3);
  assign _zz_when_ArraySlice_l166_267_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_267_3 = {1'd0, _zz_when_ArraySlice_l166_267_4};
  assign _zz__zz_when_ArraySlice_l112_267 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_267 = (_zz_when_ArraySlice_l113_267_1 - _zz_when_ArraySlice_l113_267_4);
  assign _zz_when_ArraySlice_l113_267_1 = (_zz_when_ArraySlice_l113_267_2 + _zz_when_ArraySlice_l113_267_3);
  assign _zz_when_ArraySlice_l113_267_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_267_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_267_4 = {1'd0, _zz_when_ArraySlice_l112_267};
  assign _zz__zz_when_ArraySlice_l173_267 = (_zz__zz_when_ArraySlice_l173_267_1 + _zz__zz_when_ArraySlice_l173_267_2);
  assign _zz__zz_when_ArraySlice_l173_267_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_267_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_267_3 = {1'd0, _zz_when_ArraySlice_l112_267};
  assign _zz_when_ArraySlice_l118_267_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_267 = _zz_when_ArraySlice_l118_267_1[5:0];
  assign _zz_when_ArraySlice_l173_267_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_267_1 = {1'd0, _zz_when_ArraySlice_l173_267_2};
  assign _zz_when_ArraySlice_l173_267_3 = (_zz_when_ArraySlice_l173_267_4 + _zz_when_ArraySlice_l173_267_9);
  assign _zz_when_ArraySlice_l173_267_4 = (_zz_when_ArraySlice_l173_267 - _zz_when_ArraySlice_l173_267_5);
  assign _zz_when_ArraySlice_l173_267_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_267_7);
  assign _zz_when_ArraySlice_l173_267_5 = {1'd0, _zz_when_ArraySlice_l173_267_6};
  assign _zz_when_ArraySlice_l173_267_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_267_7 = {1'd0, _zz_when_ArraySlice_l173_267_8};
  assign _zz_when_ArraySlice_l173_267_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_268 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_268_1);
  assign _zz_when_ArraySlice_l165_268_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_268 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_268_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_268_2);
  assign _zz_when_ArraySlice_l166_268_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_268_3);
  assign _zz_when_ArraySlice_l166_268_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_268 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_268 = (_zz_when_ArraySlice_l113_268_1 - _zz_when_ArraySlice_l113_268_4);
  assign _zz_when_ArraySlice_l113_268_1 = (_zz_when_ArraySlice_l113_268_2 + _zz_when_ArraySlice_l113_268_3);
  assign _zz_when_ArraySlice_l113_268_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_268_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_268_4 = {1'd0, _zz_when_ArraySlice_l112_268};
  assign _zz__zz_when_ArraySlice_l173_268 = (_zz__zz_when_ArraySlice_l173_268_1 + _zz__zz_when_ArraySlice_l173_268_2);
  assign _zz__zz_when_ArraySlice_l173_268_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_268_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_268_3 = {1'd0, _zz_when_ArraySlice_l112_268};
  assign _zz_when_ArraySlice_l118_268_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_268 = _zz_when_ArraySlice_l118_268_1[5:0];
  assign _zz_when_ArraySlice_l173_268_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_268_1 = {1'd0, _zz_when_ArraySlice_l173_268_2};
  assign _zz_when_ArraySlice_l173_268_3 = (_zz_when_ArraySlice_l173_268_4 + _zz_when_ArraySlice_l173_268_8);
  assign _zz_when_ArraySlice_l173_268_4 = (_zz_when_ArraySlice_l173_268 - _zz_when_ArraySlice_l173_268_5);
  assign _zz_when_ArraySlice_l173_268_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_268_7);
  assign _zz_when_ArraySlice_l173_268_5 = {1'd0, _zz_when_ArraySlice_l173_268_6};
  assign _zz_when_ArraySlice_l173_268_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_268_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_269 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_269_1);
  assign _zz_when_ArraySlice_l165_269_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_269_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_269 = {1'd0, _zz_when_ArraySlice_l166_269_1};
  assign _zz_when_ArraySlice_l166_269_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_269_3);
  assign _zz_when_ArraySlice_l166_269_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_269_4);
  assign _zz_when_ArraySlice_l166_269_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_269 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_269 = (_zz_when_ArraySlice_l113_269_1 - _zz_when_ArraySlice_l113_269_4);
  assign _zz_when_ArraySlice_l113_269_1 = (_zz_when_ArraySlice_l113_269_2 + _zz_when_ArraySlice_l113_269_3);
  assign _zz_when_ArraySlice_l113_269_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_269_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_269_4 = {1'd0, _zz_when_ArraySlice_l112_269};
  assign _zz__zz_when_ArraySlice_l173_269 = (_zz__zz_when_ArraySlice_l173_269_1 + _zz__zz_when_ArraySlice_l173_269_2);
  assign _zz__zz_when_ArraySlice_l173_269_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_269_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_269_3 = {1'd0, _zz_when_ArraySlice_l112_269};
  assign _zz_when_ArraySlice_l118_269_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_269 = _zz_when_ArraySlice_l118_269_1[5:0];
  assign _zz_when_ArraySlice_l173_269_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_269_1 = {2'd0, _zz_when_ArraySlice_l173_269_2};
  assign _zz_when_ArraySlice_l173_269_3 = (_zz_when_ArraySlice_l173_269_4 + _zz_when_ArraySlice_l173_269_8);
  assign _zz_when_ArraySlice_l173_269_4 = (_zz_when_ArraySlice_l173_269 - _zz_when_ArraySlice_l173_269_5);
  assign _zz_when_ArraySlice_l173_269_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_269_7);
  assign _zz_when_ArraySlice_l173_269_5 = {1'd0, _zz_when_ArraySlice_l173_269_6};
  assign _zz_when_ArraySlice_l173_269_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_269_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_270 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_270_1);
  assign _zz_when_ArraySlice_l165_270_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_270_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_270 = {1'd0, _zz_when_ArraySlice_l166_270_1};
  assign _zz_when_ArraySlice_l166_270_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_270_3);
  assign _zz_when_ArraySlice_l166_270_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_270_4);
  assign _zz_when_ArraySlice_l166_270_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_270 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_270 = (_zz_when_ArraySlice_l113_270_1 - _zz_when_ArraySlice_l113_270_4);
  assign _zz_when_ArraySlice_l113_270_1 = (_zz_when_ArraySlice_l113_270_2 + _zz_when_ArraySlice_l113_270_3);
  assign _zz_when_ArraySlice_l113_270_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_270_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_270_4 = {1'd0, _zz_when_ArraySlice_l112_270};
  assign _zz__zz_when_ArraySlice_l173_270 = (_zz__zz_when_ArraySlice_l173_270_1 + _zz__zz_when_ArraySlice_l173_270_2);
  assign _zz__zz_when_ArraySlice_l173_270_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_270_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_270_3 = {1'd0, _zz_when_ArraySlice_l112_270};
  assign _zz_when_ArraySlice_l118_270_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_270 = _zz_when_ArraySlice_l118_270_1[5:0];
  assign _zz_when_ArraySlice_l173_270_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_270_1 = {2'd0, _zz_when_ArraySlice_l173_270_2};
  assign _zz_when_ArraySlice_l173_270_3 = (_zz_when_ArraySlice_l173_270_4 + _zz_when_ArraySlice_l173_270_8);
  assign _zz_when_ArraySlice_l173_270_4 = (_zz_when_ArraySlice_l173_270 - _zz_when_ArraySlice_l173_270_5);
  assign _zz_when_ArraySlice_l173_270_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_270_7);
  assign _zz_when_ArraySlice_l173_270_5 = {1'd0, _zz_when_ArraySlice_l173_270_6};
  assign _zz_when_ArraySlice_l173_270_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_270_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_271 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_271_1);
  assign _zz_when_ArraySlice_l165_271_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_271_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_271 = {2'd0, _zz_when_ArraySlice_l166_271_1};
  assign _zz_when_ArraySlice_l166_271_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_271_3);
  assign _zz_when_ArraySlice_l166_271_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_271_4);
  assign _zz_when_ArraySlice_l166_271_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_271 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_271 = (_zz_when_ArraySlice_l113_271_1 - _zz_when_ArraySlice_l113_271_4);
  assign _zz_when_ArraySlice_l113_271_1 = (_zz_when_ArraySlice_l113_271_2 + _zz_when_ArraySlice_l113_271_3);
  assign _zz_when_ArraySlice_l113_271_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_271_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_271_4 = {1'd0, _zz_when_ArraySlice_l112_271};
  assign _zz__zz_when_ArraySlice_l173_271 = (_zz__zz_when_ArraySlice_l173_271_1 + _zz__zz_when_ArraySlice_l173_271_2);
  assign _zz__zz_when_ArraySlice_l173_271_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_271_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_271_3 = {1'd0, _zz_when_ArraySlice_l112_271};
  assign _zz_when_ArraySlice_l118_271_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_271 = _zz_when_ArraySlice_l118_271_1[5:0];
  assign _zz_when_ArraySlice_l173_271_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_271_1 = {3'd0, _zz_when_ArraySlice_l173_271_2};
  assign _zz_when_ArraySlice_l173_271_3 = (_zz_when_ArraySlice_l173_271_4 + _zz_when_ArraySlice_l173_271_8);
  assign _zz_when_ArraySlice_l173_271_4 = (_zz_when_ArraySlice_l173_271 - _zz_when_ArraySlice_l173_271_5);
  assign _zz_when_ArraySlice_l173_271_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_271_7);
  assign _zz_when_ArraySlice_l173_271_5 = {1'd0, _zz_when_ArraySlice_l173_271_6};
  assign _zz_when_ArraySlice_l173_271_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_271_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l288_2_1 = (_zz_when_ArraySlice_l288_2_2 + _zz_when_ArraySlice_l288_2_7);
  assign _zz_when_ArraySlice_l288_2_2 = (_zz_when_ArraySlice_l288_2_3 + _zz_when_ArraySlice_l288_2_5);
  assign _zz_when_ArraySlice_l288_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l288_2_4);
  assign _zz_when_ArraySlice_l288_2_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l288_2_5 = {5'd0, _zz_when_ArraySlice_l288_2_6};
  assign _zz_when_ArraySlice_l288_2_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l288_2_7 = {1'd0, _zz_when_ArraySlice_l288_2_8};
  assign _zz_selectReadFifo_2_57 = 1'b1;
  assign _zz_selectReadFifo_2_56 = {5'd0, _zz_selectReadFifo_2_57};
  assign _zz_when_ArraySlice_l292_2_1 = (_zz_when_ArraySlice_l292_2_2 % aReg);
  assign _zz_when_ArraySlice_l292_2_2 = (handshakeTimes_2_value + _zz_when_ArraySlice_l292_2_3);
  assign _zz_when_ArraySlice_l292_2_4 = 1'b1;
  assign _zz_when_ArraySlice_l292_2_3 = {12'd0, _zz_when_ArraySlice_l292_2_4};
  assign _zz_when_ArraySlice_l303_2_2 = (_zz_when_ArraySlice_l303_2_3 - _zz_when_ArraySlice_l303_2_4);
  assign _zz_when_ArraySlice_l303_2_1 = {7'd0, _zz_when_ArraySlice_l303_2_2};
  assign _zz_when_ArraySlice_l303_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l303_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l303_2_4 = {5'd0, _zz_when_ArraySlice_l303_2_5};
  assign _zz__zz_when_ArraySlice_l94_32 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_32 = (_zz_when_ArraySlice_l95_32_1 - _zz_when_ArraySlice_l95_32_4);
  assign _zz_when_ArraySlice_l95_32_1 = (_zz_when_ArraySlice_l95_32_2 + _zz_when_ArraySlice_l95_32_3);
  assign _zz_when_ArraySlice_l95_32_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_32_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_32_4 = {1'd0, _zz_when_ArraySlice_l94_32};
  assign _zz__zz_when_ArraySlice_l304_2_1 = (_zz__zz_when_ArraySlice_l304_2_2 + _zz__zz_when_ArraySlice_l304_2_3);
  assign _zz__zz_when_ArraySlice_l304_2_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l304_2_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l304_2_4 = {1'd0, _zz_when_ArraySlice_l94_32};
  assign _zz_when_ArraySlice_l99_32_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_32 = _zz_when_ArraySlice_l99_32_1[5:0];
  assign _zz_when_ArraySlice_l304_2_1 = (outSliceNumb_2_value + _zz_when_ArraySlice_l304_2_2);
  assign _zz_when_ArraySlice_l304_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l304_2_2 = {6'd0, _zz_when_ArraySlice_l304_2_3};
  assign _zz_when_ArraySlice_l304_2_4 = (_zz_when_ArraySlice_l304_2 / aReg);
  assign _zz_selectReadFifo_2_58 = (selectReadFifo_2 - _zz_selectReadFifo_2_59);
  assign _zz_selectReadFifo_2_59 = {3'd0, bReg};
  assign _zz_selectReadFifo_2_61 = 1'b1;
  assign _zz_selectReadFifo_2_60 = {5'd0, _zz_selectReadFifo_2_61};
  assign _zz_when_ArraySlice_l165_272 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_272_1);
  assign _zz_when_ArraySlice_l165_272_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_272_1 = {3'd0, _zz_when_ArraySlice_l165_272_2};
  assign _zz_when_ArraySlice_l166_272 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_272_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_272_3);
  assign _zz_when_ArraySlice_l166_272_1 = {1'd0, _zz_when_ArraySlice_l166_272_2};
  assign _zz_when_ArraySlice_l166_272_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_272_4);
  assign _zz_when_ArraySlice_l166_272_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_272_4 = {3'd0, _zz_when_ArraySlice_l166_272_5};
  assign _zz__zz_when_ArraySlice_l112_272 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_272 = (_zz_when_ArraySlice_l113_272_1 - _zz_when_ArraySlice_l113_272_4);
  assign _zz_when_ArraySlice_l113_272_1 = (_zz_when_ArraySlice_l113_272_2 + _zz_when_ArraySlice_l113_272_3);
  assign _zz_when_ArraySlice_l113_272_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_272_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_272_4 = {1'd0, _zz_when_ArraySlice_l112_272};
  assign _zz__zz_when_ArraySlice_l173_272 = (_zz__zz_when_ArraySlice_l173_272_1 + _zz__zz_when_ArraySlice_l173_272_2);
  assign _zz__zz_when_ArraySlice_l173_272_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_272_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_272_3 = {1'd0, _zz_when_ArraySlice_l112_272};
  assign _zz_when_ArraySlice_l118_272_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_272 = _zz_when_ArraySlice_l118_272_1[5:0];
  assign _zz_when_ArraySlice_l173_272_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_272_2 = (_zz_when_ArraySlice_l173_272_3 + _zz_when_ArraySlice_l173_272_8);
  assign _zz_when_ArraySlice_l173_272_3 = (_zz_when_ArraySlice_l173_272 - _zz_when_ArraySlice_l173_272_4);
  assign _zz_when_ArraySlice_l173_272_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_272_6);
  assign _zz_when_ArraySlice_l173_272_4 = {1'd0, _zz_when_ArraySlice_l173_272_5};
  assign _zz_when_ArraySlice_l173_272_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_272_6 = {3'd0, _zz_when_ArraySlice_l173_272_7};
  assign _zz_when_ArraySlice_l173_272_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_273 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_273_1);
  assign _zz_when_ArraySlice_l165_273_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_273_1 = {2'd0, _zz_when_ArraySlice_l165_273_2};
  assign _zz_when_ArraySlice_l166_273 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_273_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_273_2);
  assign _zz_when_ArraySlice_l166_273_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_273_3);
  assign _zz_when_ArraySlice_l166_273_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_273_3 = {2'd0, _zz_when_ArraySlice_l166_273_4};
  assign _zz__zz_when_ArraySlice_l112_273 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_273 = (_zz_when_ArraySlice_l113_273_1 - _zz_when_ArraySlice_l113_273_4);
  assign _zz_when_ArraySlice_l113_273_1 = (_zz_when_ArraySlice_l113_273_2 + _zz_when_ArraySlice_l113_273_3);
  assign _zz_when_ArraySlice_l113_273_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_273_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_273_4 = {1'd0, _zz_when_ArraySlice_l112_273};
  assign _zz__zz_when_ArraySlice_l173_273 = (_zz__zz_when_ArraySlice_l173_273_1 + _zz__zz_when_ArraySlice_l173_273_2);
  assign _zz__zz_when_ArraySlice_l173_273_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_273_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_273_3 = {1'd0, _zz_when_ArraySlice_l112_273};
  assign _zz_when_ArraySlice_l118_273_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_273 = _zz_when_ArraySlice_l118_273_1[5:0];
  assign _zz_when_ArraySlice_l173_273_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_273_1 = {1'd0, _zz_when_ArraySlice_l173_273_2};
  assign _zz_when_ArraySlice_l173_273_3 = (_zz_when_ArraySlice_l173_273_4 + _zz_when_ArraySlice_l173_273_9);
  assign _zz_when_ArraySlice_l173_273_4 = (_zz_when_ArraySlice_l173_273 - _zz_when_ArraySlice_l173_273_5);
  assign _zz_when_ArraySlice_l173_273_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_273_7);
  assign _zz_when_ArraySlice_l173_273_5 = {1'd0, _zz_when_ArraySlice_l173_273_6};
  assign _zz_when_ArraySlice_l173_273_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_273_7 = {2'd0, _zz_when_ArraySlice_l173_273_8};
  assign _zz_when_ArraySlice_l173_273_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_274 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_274_1);
  assign _zz_when_ArraySlice_l165_274_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_274_1 = {1'd0, _zz_when_ArraySlice_l165_274_2};
  assign _zz_when_ArraySlice_l166_274 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_274_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_274_2);
  assign _zz_when_ArraySlice_l166_274_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_274_3);
  assign _zz_when_ArraySlice_l166_274_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_274_3 = {1'd0, _zz_when_ArraySlice_l166_274_4};
  assign _zz__zz_when_ArraySlice_l112_274 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_274 = (_zz_when_ArraySlice_l113_274_1 - _zz_when_ArraySlice_l113_274_4);
  assign _zz_when_ArraySlice_l113_274_1 = (_zz_when_ArraySlice_l113_274_2 + _zz_when_ArraySlice_l113_274_3);
  assign _zz_when_ArraySlice_l113_274_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_274_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_274_4 = {1'd0, _zz_when_ArraySlice_l112_274};
  assign _zz__zz_when_ArraySlice_l173_274 = (_zz__zz_when_ArraySlice_l173_274_1 + _zz__zz_when_ArraySlice_l173_274_2);
  assign _zz__zz_when_ArraySlice_l173_274_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_274_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_274_3 = {1'd0, _zz_when_ArraySlice_l112_274};
  assign _zz_when_ArraySlice_l118_274_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_274 = _zz_when_ArraySlice_l118_274_1[5:0];
  assign _zz_when_ArraySlice_l173_274_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_274_1 = {1'd0, _zz_when_ArraySlice_l173_274_2};
  assign _zz_when_ArraySlice_l173_274_3 = (_zz_when_ArraySlice_l173_274_4 + _zz_when_ArraySlice_l173_274_9);
  assign _zz_when_ArraySlice_l173_274_4 = (_zz_when_ArraySlice_l173_274 - _zz_when_ArraySlice_l173_274_5);
  assign _zz_when_ArraySlice_l173_274_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_274_7);
  assign _zz_when_ArraySlice_l173_274_5 = {1'd0, _zz_when_ArraySlice_l173_274_6};
  assign _zz_when_ArraySlice_l173_274_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_274_7 = {1'd0, _zz_when_ArraySlice_l173_274_8};
  assign _zz_when_ArraySlice_l173_274_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_275 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_275_1);
  assign _zz_when_ArraySlice_l165_275_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_275_1 = {1'd0, _zz_when_ArraySlice_l165_275_2};
  assign _zz_when_ArraySlice_l166_275 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_275_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_275_2);
  assign _zz_when_ArraySlice_l166_275_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_275_3);
  assign _zz_when_ArraySlice_l166_275_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_275_3 = {1'd0, _zz_when_ArraySlice_l166_275_4};
  assign _zz__zz_when_ArraySlice_l112_275 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_275 = (_zz_when_ArraySlice_l113_275_1 - _zz_when_ArraySlice_l113_275_4);
  assign _zz_when_ArraySlice_l113_275_1 = (_zz_when_ArraySlice_l113_275_2 + _zz_when_ArraySlice_l113_275_3);
  assign _zz_when_ArraySlice_l113_275_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_275_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_275_4 = {1'd0, _zz_when_ArraySlice_l112_275};
  assign _zz__zz_when_ArraySlice_l173_275 = (_zz__zz_when_ArraySlice_l173_275_1 + _zz__zz_when_ArraySlice_l173_275_2);
  assign _zz__zz_when_ArraySlice_l173_275_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_275_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_275_3 = {1'd0, _zz_when_ArraySlice_l112_275};
  assign _zz_when_ArraySlice_l118_275_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_275 = _zz_when_ArraySlice_l118_275_1[5:0];
  assign _zz_when_ArraySlice_l173_275_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_275_1 = {1'd0, _zz_when_ArraySlice_l173_275_2};
  assign _zz_when_ArraySlice_l173_275_3 = (_zz_when_ArraySlice_l173_275_4 + _zz_when_ArraySlice_l173_275_9);
  assign _zz_when_ArraySlice_l173_275_4 = (_zz_when_ArraySlice_l173_275 - _zz_when_ArraySlice_l173_275_5);
  assign _zz_when_ArraySlice_l173_275_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_275_7);
  assign _zz_when_ArraySlice_l173_275_5 = {1'd0, _zz_when_ArraySlice_l173_275_6};
  assign _zz_when_ArraySlice_l173_275_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_275_7 = {1'd0, _zz_when_ArraySlice_l173_275_8};
  assign _zz_when_ArraySlice_l173_275_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_276 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_276_1);
  assign _zz_when_ArraySlice_l165_276_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_276 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_276_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_276_2);
  assign _zz_when_ArraySlice_l166_276_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_276_3);
  assign _zz_when_ArraySlice_l166_276_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_276 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_276 = (_zz_when_ArraySlice_l113_276_1 - _zz_when_ArraySlice_l113_276_4);
  assign _zz_when_ArraySlice_l113_276_1 = (_zz_when_ArraySlice_l113_276_2 + _zz_when_ArraySlice_l113_276_3);
  assign _zz_when_ArraySlice_l113_276_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_276_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_276_4 = {1'd0, _zz_when_ArraySlice_l112_276};
  assign _zz__zz_when_ArraySlice_l173_276 = (_zz__zz_when_ArraySlice_l173_276_1 + _zz__zz_when_ArraySlice_l173_276_2);
  assign _zz__zz_when_ArraySlice_l173_276_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_276_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_276_3 = {1'd0, _zz_when_ArraySlice_l112_276};
  assign _zz_when_ArraySlice_l118_276_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_276 = _zz_when_ArraySlice_l118_276_1[5:0];
  assign _zz_when_ArraySlice_l173_276_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_276_1 = {1'd0, _zz_when_ArraySlice_l173_276_2};
  assign _zz_when_ArraySlice_l173_276_3 = (_zz_when_ArraySlice_l173_276_4 + _zz_when_ArraySlice_l173_276_8);
  assign _zz_when_ArraySlice_l173_276_4 = (_zz_when_ArraySlice_l173_276 - _zz_when_ArraySlice_l173_276_5);
  assign _zz_when_ArraySlice_l173_276_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_276_7);
  assign _zz_when_ArraySlice_l173_276_5 = {1'd0, _zz_when_ArraySlice_l173_276_6};
  assign _zz_when_ArraySlice_l173_276_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_276_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_277 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_277_1);
  assign _zz_when_ArraySlice_l165_277_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_277_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_277 = {1'd0, _zz_when_ArraySlice_l166_277_1};
  assign _zz_when_ArraySlice_l166_277_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_277_3);
  assign _zz_when_ArraySlice_l166_277_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_277_4);
  assign _zz_when_ArraySlice_l166_277_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_277 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_277 = (_zz_when_ArraySlice_l113_277_1 - _zz_when_ArraySlice_l113_277_4);
  assign _zz_when_ArraySlice_l113_277_1 = (_zz_when_ArraySlice_l113_277_2 + _zz_when_ArraySlice_l113_277_3);
  assign _zz_when_ArraySlice_l113_277_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_277_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_277_4 = {1'd0, _zz_when_ArraySlice_l112_277};
  assign _zz__zz_when_ArraySlice_l173_277 = (_zz__zz_when_ArraySlice_l173_277_1 + _zz__zz_when_ArraySlice_l173_277_2);
  assign _zz__zz_when_ArraySlice_l173_277_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_277_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_277_3 = {1'd0, _zz_when_ArraySlice_l112_277};
  assign _zz_when_ArraySlice_l118_277_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_277 = _zz_when_ArraySlice_l118_277_1[5:0];
  assign _zz_when_ArraySlice_l173_277_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_277_1 = {2'd0, _zz_when_ArraySlice_l173_277_2};
  assign _zz_when_ArraySlice_l173_277_3 = (_zz_when_ArraySlice_l173_277_4 + _zz_when_ArraySlice_l173_277_8);
  assign _zz_when_ArraySlice_l173_277_4 = (_zz_when_ArraySlice_l173_277 - _zz_when_ArraySlice_l173_277_5);
  assign _zz_when_ArraySlice_l173_277_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_277_7);
  assign _zz_when_ArraySlice_l173_277_5 = {1'd0, _zz_when_ArraySlice_l173_277_6};
  assign _zz_when_ArraySlice_l173_277_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_277_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_278 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_278_1);
  assign _zz_when_ArraySlice_l165_278_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_278_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_278 = {1'd0, _zz_when_ArraySlice_l166_278_1};
  assign _zz_when_ArraySlice_l166_278_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_278_3);
  assign _zz_when_ArraySlice_l166_278_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_278_4);
  assign _zz_when_ArraySlice_l166_278_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_278 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_278 = (_zz_when_ArraySlice_l113_278_1 - _zz_when_ArraySlice_l113_278_4);
  assign _zz_when_ArraySlice_l113_278_1 = (_zz_when_ArraySlice_l113_278_2 + _zz_when_ArraySlice_l113_278_3);
  assign _zz_when_ArraySlice_l113_278_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_278_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_278_4 = {1'd0, _zz_when_ArraySlice_l112_278};
  assign _zz__zz_when_ArraySlice_l173_278 = (_zz__zz_when_ArraySlice_l173_278_1 + _zz__zz_when_ArraySlice_l173_278_2);
  assign _zz__zz_when_ArraySlice_l173_278_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_278_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_278_3 = {1'd0, _zz_when_ArraySlice_l112_278};
  assign _zz_when_ArraySlice_l118_278_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_278 = _zz_when_ArraySlice_l118_278_1[5:0];
  assign _zz_when_ArraySlice_l173_278_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_278_1 = {2'd0, _zz_when_ArraySlice_l173_278_2};
  assign _zz_when_ArraySlice_l173_278_3 = (_zz_when_ArraySlice_l173_278_4 + _zz_when_ArraySlice_l173_278_8);
  assign _zz_when_ArraySlice_l173_278_4 = (_zz_when_ArraySlice_l173_278 - _zz_when_ArraySlice_l173_278_5);
  assign _zz_when_ArraySlice_l173_278_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_278_7);
  assign _zz_when_ArraySlice_l173_278_5 = {1'd0, _zz_when_ArraySlice_l173_278_6};
  assign _zz_when_ArraySlice_l173_278_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_278_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_279 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_279_1);
  assign _zz_when_ArraySlice_l165_279_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_279_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_279 = {2'd0, _zz_when_ArraySlice_l166_279_1};
  assign _zz_when_ArraySlice_l166_279_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_279_3);
  assign _zz_when_ArraySlice_l166_279_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_279_4);
  assign _zz_when_ArraySlice_l166_279_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_279 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_279 = (_zz_when_ArraySlice_l113_279_1 - _zz_when_ArraySlice_l113_279_4);
  assign _zz_when_ArraySlice_l113_279_1 = (_zz_when_ArraySlice_l113_279_2 + _zz_when_ArraySlice_l113_279_3);
  assign _zz_when_ArraySlice_l113_279_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_279_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_279_4 = {1'd0, _zz_when_ArraySlice_l112_279};
  assign _zz__zz_when_ArraySlice_l173_279 = (_zz__zz_when_ArraySlice_l173_279_1 + _zz__zz_when_ArraySlice_l173_279_2);
  assign _zz__zz_when_ArraySlice_l173_279_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_279_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_279_3 = {1'd0, _zz_when_ArraySlice_l112_279};
  assign _zz_when_ArraySlice_l118_279_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_279 = _zz_when_ArraySlice_l118_279_1[5:0];
  assign _zz_when_ArraySlice_l173_279_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_279_1 = {3'd0, _zz_when_ArraySlice_l173_279_2};
  assign _zz_when_ArraySlice_l173_279_3 = (_zz_when_ArraySlice_l173_279_4 + _zz_when_ArraySlice_l173_279_8);
  assign _zz_when_ArraySlice_l173_279_4 = (_zz_when_ArraySlice_l173_279 - _zz_when_ArraySlice_l173_279_5);
  assign _zz_when_ArraySlice_l173_279_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_279_7);
  assign _zz_when_ArraySlice_l173_279_5 = {1'd0, _zz_when_ArraySlice_l173_279_6};
  assign _zz_when_ArraySlice_l173_279_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_279_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_2_63 = 1'b1;
  assign _zz_selectReadFifo_2_62 = {5'd0, _zz_selectReadFifo_2_63};
  assign _zz_when_ArraySlice_l315_2_1 = (_zz_when_ArraySlice_l315_2_2 % aReg);
  assign _zz_when_ArraySlice_l315_2_2 = (handshakeTimes_2_value + _zz_when_ArraySlice_l315_2_3);
  assign _zz_when_ArraySlice_l315_2_4 = 1'b1;
  assign _zz_when_ArraySlice_l315_2_3 = {12'd0, _zz_when_ArraySlice_l315_2_4};
  assign _zz_when_ArraySlice_l301_2_1 = (selectReadFifo_2 + _zz_when_ArraySlice_l301_2_2);
  assign _zz_when_ArraySlice_l301_2_3 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l301_2_2 = {1'd0, _zz_when_ArraySlice_l301_2_3};
  assign _zz_when_ArraySlice_l322_2_2 = (_zz_when_ArraySlice_l322_2_3 - _zz_when_ArraySlice_l322_2_4);
  assign _zz_when_ArraySlice_l322_2_1 = {7'd0, _zz_when_ArraySlice_l322_2_2};
  assign _zz_when_ArraySlice_l322_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l322_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l322_2_4 = {5'd0, _zz_when_ArraySlice_l322_2_5};
  assign _zz_when_ArraySlice_l240_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l240_3_1);
  assign _zz_when_ArraySlice_l240_3_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l240_3_1 = {1'd0, _zz_when_ArraySlice_l240_3_2};
  assign _zz_when_ArraySlice_l241_3_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l241_3_3);
  assign _zz_when_ArraySlice_l241_3_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l241_3_3 = {1'd0, _zz_when_ArraySlice_l241_3_4};
  assign _zz__zz_outputStreamArrayData_3_valid_1_2 = (bReg * 2'b11);
  assign _zz__zz_outputStreamArrayData_3_valid_1_1 = {1'd0, _zz__zz_outputStreamArrayData_3_valid_1_2};
  assign _zz_when_ArraySlice_l247_3_2 = 1'b1;
  assign _zz_when_ArraySlice_l247_3_1 = {6'd0, _zz_when_ArraySlice_l247_3_2};
  assign _zz_when_ArraySlice_l247_3_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l247_3_5);
  assign _zz_when_ArraySlice_l247_3_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l247_3_5 = {1'd0, _zz_when_ArraySlice_l247_3_6};
  assign _zz_when_ArraySlice_l248_3_2 = (_zz_when_ArraySlice_l248_3_3 - _zz_when_ArraySlice_l248_3_4);
  assign _zz_when_ArraySlice_l248_3_1 = {7'd0, _zz_when_ArraySlice_l248_3_2};
  assign _zz_when_ArraySlice_l248_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l248_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l248_3_4 = {5'd0, _zz_when_ArraySlice_l248_3_5};
  assign _zz_selectReadFifo_3_32 = (selectReadFifo_3 - _zz_selectReadFifo_3_33);
  assign _zz_selectReadFifo_3_33 = {3'd0, bReg};
  assign _zz_selectReadFifo_3_35 = 1'b1;
  assign _zz_selectReadFifo_3_34 = {5'd0, _zz_selectReadFifo_3_35};
  assign _zz_selectReadFifo_3_37 = 1'b1;
  assign _zz_selectReadFifo_3_36 = {5'd0, _zz_selectReadFifo_3_37};
  assign _zz_when_ArraySlice_l251_3_1 = (_zz_when_ArraySlice_l251_3_2 % aReg);
  assign _zz_when_ArraySlice_l251_3_2 = (handshakeTimes_3_value + _zz_when_ArraySlice_l251_3_3);
  assign _zz_when_ArraySlice_l251_3_4 = 1'b1;
  assign _zz_when_ArraySlice_l251_3_3 = {12'd0, _zz_when_ArraySlice_l251_3_4};
  assign _zz_when_ArraySlice_l256_3_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l256_3_3);
  assign _zz_when_ArraySlice_l256_3_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l256_3_3 = {1'd0, _zz_when_ArraySlice_l256_3_4};
  assign _zz_when_ArraySlice_l256_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l256_3_5 = {6'd0, _zz_when_ArraySlice_l256_3_6};
  assign _zz_when_ArraySlice_l257_3_2 = (_zz_when_ArraySlice_l257_3_3 - _zz_when_ArraySlice_l257_3_4);
  assign _zz_when_ArraySlice_l257_3_1 = {7'd0, _zz_when_ArraySlice_l257_3_2};
  assign _zz_when_ArraySlice_l257_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l257_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l257_3_4 = {5'd0, _zz_when_ArraySlice_l257_3_5};
  assign _zz__zz_when_ArraySlice_l94_33 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_33 = (_zz_when_ArraySlice_l95_33_1 - _zz_when_ArraySlice_l95_33_4);
  assign _zz_when_ArraySlice_l95_33_1 = (_zz_when_ArraySlice_l95_33_2 + _zz_when_ArraySlice_l95_33_3);
  assign _zz_when_ArraySlice_l95_33_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_33_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_33_4 = {1'd0, _zz_when_ArraySlice_l94_33};
  assign _zz__zz_when_ArraySlice_l259_3_1 = (_zz__zz_when_ArraySlice_l259_3_2 + _zz__zz_when_ArraySlice_l259_3_3);
  assign _zz__zz_when_ArraySlice_l259_3_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l259_3_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l259_3_4 = {1'd0, _zz_when_ArraySlice_l94_33};
  assign _zz_when_ArraySlice_l99_33_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_33 = _zz_when_ArraySlice_l99_33_1[5:0];
  assign _zz_when_ArraySlice_l259_3_1 = (outSliceNumb_3_value + _zz_when_ArraySlice_l259_3_2);
  assign _zz_when_ArraySlice_l259_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l259_3_2 = {6'd0, _zz_when_ArraySlice_l259_3_3};
  assign _zz_when_ArraySlice_l259_3_4 = (_zz_when_ArraySlice_l259_3 / aReg);
  assign _zz_selectReadFifo_3_38 = (selectReadFifo_3 - _zz_selectReadFifo_3_39);
  assign _zz_selectReadFifo_3_39 = {3'd0, bReg};
  assign _zz_selectReadFifo_3_41 = 1'b1;
  assign _zz_selectReadFifo_3_40 = {5'd0, _zz_selectReadFifo_3_41};
  assign _zz_selectReadFifo_3_42 = (selectReadFifo_3 + _zz_selectReadFifo_3_43);
  assign _zz_selectReadFifo_3_43 = (3'b111 * bReg);
  assign _zz_selectReadFifo_3_45 = 1'b1;
  assign _zz_selectReadFifo_3_44 = {5'd0, _zz_selectReadFifo_3_45};
  assign _zz_when_ArraySlice_l165_280 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_280_1);
  assign _zz_when_ArraySlice_l165_280_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_280_1 = {3'd0, _zz_when_ArraySlice_l165_280_2};
  assign _zz_when_ArraySlice_l166_280 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_280_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_280_3);
  assign _zz_when_ArraySlice_l166_280_1 = {1'd0, _zz_when_ArraySlice_l166_280_2};
  assign _zz_when_ArraySlice_l166_280_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_280_4);
  assign _zz_when_ArraySlice_l166_280_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_280_4 = {3'd0, _zz_when_ArraySlice_l166_280_5};
  assign _zz__zz_when_ArraySlice_l112_280 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_280 = (_zz_when_ArraySlice_l113_280_1 - _zz_when_ArraySlice_l113_280_4);
  assign _zz_when_ArraySlice_l113_280_1 = (_zz_when_ArraySlice_l113_280_2 + _zz_when_ArraySlice_l113_280_3);
  assign _zz_when_ArraySlice_l113_280_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_280_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_280_4 = {1'd0, _zz_when_ArraySlice_l112_280};
  assign _zz__zz_when_ArraySlice_l173_280 = (_zz__zz_when_ArraySlice_l173_280_1 + _zz__zz_when_ArraySlice_l173_280_2);
  assign _zz__zz_when_ArraySlice_l173_280_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_280_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_280_3 = {1'd0, _zz_when_ArraySlice_l112_280};
  assign _zz_when_ArraySlice_l118_280_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_280 = _zz_when_ArraySlice_l118_280_1[5:0];
  assign _zz_when_ArraySlice_l173_280_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_280_2 = (_zz_when_ArraySlice_l173_280_3 + _zz_when_ArraySlice_l173_280_8);
  assign _zz_when_ArraySlice_l173_280_3 = (_zz_when_ArraySlice_l173_280 - _zz_when_ArraySlice_l173_280_4);
  assign _zz_when_ArraySlice_l173_280_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_280_6);
  assign _zz_when_ArraySlice_l173_280_4 = {1'd0, _zz_when_ArraySlice_l173_280_5};
  assign _zz_when_ArraySlice_l173_280_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_280_6 = {3'd0, _zz_when_ArraySlice_l173_280_7};
  assign _zz_when_ArraySlice_l173_280_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_281 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_281_1);
  assign _zz_when_ArraySlice_l165_281_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_281_1 = {2'd0, _zz_when_ArraySlice_l165_281_2};
  assign _zz_when_ArraySlice_l166_281 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_281_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_281_2);
  assign _zz_when_ArraySlice_l166_281_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_281_3);
  assign _zz_when_ArraySlice_l166_281_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_281_3 = {2'd0, _zz_when_ArraySlice_l166_281_4};
  assign _zz__zz_when_ArraySlice_l112_281 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_281 = (_zz_when_ArraySlice_l113_281_1 - _zz_when_ArraySlice_l113_281_4);
  assign _zz_when_ArraySlice_l113_281_1 = (_zz_when_ArraySlice_l113_281_2 + _zz_when_ArraySlice_l113_281_3);
  assign _zz_when_ArraySlice_l113_281_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_281_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_281_4 = {1'd0, _zz_when_ArraySlice_l112_281};
  assign _zz__zz_when_ArraySlice_l173_281 = (_zz__zz_when_ArraySlice_l173_281_1 + _zz__zz_when_ArraySlice_l173_281_2);
  assign _zz__zz_when_ArraySlice_l173_281_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_281_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_281_3 = {1'd0, _zz_when_ArraySlice_l112_281};
  assign _zz_when_ArraySlice_l118_281_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_281 = _zz_when_ArraySlice_l118_281_1[5:0];
  assign _zz_when_ArraySlice_l173_281_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_281_1 = {1'd0, _zz_when_ArraySlice_l173_281_2};
  assign _zz_when_ArraySlice_l173_281_3 = (_zz_when_ArraySlice_l173_281_4 + _zz_when_ArraySlice_l173_281_9);
  assign _zz_when_ArraySlice_l173_281_4 = (_zz_when_ArraySlice_l173_281 - _zz_when_ArraySlice_l173_281_5);
  assign _zz_when_ArraySlice_l173_281_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_281_7);
  assign _zz_when_ArraySlice_l173_281_5 = {1'd0, _zz_when_ArraySlice_l173_281_6};
  assign _zz_when_ArraySlice_l173_281_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_281_7 = {2'd0, _zz_when_ArraySlice_l173_281_8};
  assign _zz_when_ArraySlice_l173_281_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_282 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_282_1);
  assign _zz_when_ArraySlice_l165_282_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_282_1 = {1'd0, _zz_when_ArraySlice_l165_282_2};
  assign _zz_when_ArraySlice_l166_282 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_282_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_282_2);
  assign _zz_when_ArraySlice_l166_282_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_282_3);
  assign _zz_when_ArraySlice_l166_282_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_282_3 = {1'd0, _zz_when_ArraySlice_l166_282_4};
  assign _zz__zz_when_ArraySlice_l112_282 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_282 = (_zz_when_ArraySlice_l113_282_1 - _zz_when_ArraySlice_l113_282_4);
  assign _zz_when_ArraySlice_l113_282_1 = (_zz_when_ArraySlice_l113_282_2 + _zz_when_ArraySlice_l113_282_3);
  assign _zz_when_ArraySlice_l113_282_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_282_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_282_4 = {1'd0, _zz_when_ArraySlice_l112_282};
  assign _zz__zz_when_ArraySlice_l173_282 = (_zz__zz_when_ArraySlice_l173_282_1 + _zz__zz_when_ArraySlice_l173_282_2);
  assign _zz__zz_when_ArraySlice_l173_282_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_282_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_282_3 = {1'd0, _zz_when_ArraySlice_l112_282};
  assign _zz_when_ArraySlice_l118_282_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_282 = _zz_when_ArraySlice_l118_282_1[5:0];
  assign _zz_when_ArraySlice_l173_282_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_282_1 = {1'd0, _zz_when_ArraySlice_l173_282_2};
  assign _zz_when_ArraySlice_l173_282_3 = (_zz_when_ArraySlice_l173_282_4 + _zz_when_ArraySlice_l173_282_9);
  assign _zz_when_ArraySlice_l173_282_4 = (_zz_when_ArraySlice_l173_282 - _zz_when_ArraySlice_l173_282_5);
  assign _zz_when_ArraySlice_l173_282_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_282_7);
  assign _zz_when_ArraySlice_l173_282_5 = {1'd0, _zz_when_ArraySlice_l173_282_6};
  assign _zz_when_ArraySlice_l173_282_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_282_7 = {1'd0, _zz_when_ArraySlice_l173_282_8};
  assign _zz_when_ArraySlice_l173_282_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_283 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_283_1);
  assign _zz_when_ArraySlice_l165_283_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_283_1 = {1'd0, _zz_when_ArraySlice_l165_283_2};
  assign _zz_when_ArraySlice_l166_283 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_283_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_283_2);
  assign _zz_when_ArraySlice_l166_283_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_283_3);
  assign _zz_when_ArraySlice_l166_283_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_283_3 = {1'd0, _zz_when_ArraySlice_l166_283_4};
  assign _zz__zz_when_ArraySlice_l112_283 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_283 = (_zz_when_ArraySlice_l113_283_1 - _zz_when_ArraySlice_l113_283_4);
  assign _zz_when_ArraySlice_l113_283_1 = (_zz_when_ArraySlice_l113_283_2 + _zz_when_ArraySlice_l113_283_3);
  assign _zz_when_ArraySlice_l113_283_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_283_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_283_4 = {1'd0, _zz_when_ArraySlice_l112_283};
  assign _zz__zz_when_ArraySlice_l173_283 = (_zz__zz_when_ArraySlice_l173_283_1 + _zz__zz_when_ArraySlice_l173_283_2);
  assign _zz__zz_when_ArraySlice_l173_283_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_283_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_283_3 = {1'd0, _zz_when_ArraySlice_l112_283};
  assign _zz_when_ArraySlice_l118_283_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_283 = _zz_when_ArraySlice_l118_283_1[5:0];
  assign _zz_when_ArraySlice_l173_283_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_283_1 = {1'd0, _zz_when_ArraySlice_l173_283_2};
  assign _zz_when_ArraySlice_l173_283_3 = (_zz_when_ArraySlice_l173_283_4 + _zz_when_ArraySlice_l173_283_9);
  assign _zz_when_ArraySlice_l173_283_4 = (_zz_when_ArraySlice_l173_283 - _zz_when_ArraySlice_l173_283_5);
  assign _zz_when_ArraySlice_l173_283_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_283_7);
  assign _zz_when_ArraySlice_l173_283_5 = {1'd0, _zz_when_ArraySlice_l173_283_6};
  assign _zz_when_ArraySlice_l173_283_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_283_7 = {1'd0, _zz_when_ArraySlice_l173_283_8};
  assign _zz_when_ArraySlice_l173_283_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_284 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_284_1);
  assign _zz_when_ArraySlice_l165_284_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_284 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_284_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_284_2);
  assign _zz_when_ArraySlice_l166_284_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_284_3);
  assign _zz_when_ArraySlice_l166_284_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_284 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_284 = (_zz_when_ArraySlice_l113_284_1 - _zz_when_ArraySlice_l113_284_4);
  assign _zz_when_ArraySlice_l113_284_1 = (_zz_when_ArraySlice_l113_284_2 + _zz_when_ArraySlice_l113_284_3);
  assign _zz_when_ArraySlice_l113_284_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_284_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_284_4 = {1'd0, _zz_when_ArraySlice_l112_284};
  assign _zz__zz_when_ArraySlice_l173_284 = (_zz__zz_when_ArraySlice_l173_284_1 + _zz__zz_when_ArraySlice_l173_284_2);
  assign _zz__zz_when_ArraySlice_l173_284_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_284_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_284_3 = {1'd0, _zz_when_ArraySlice_l112_284};
  assign _zz_when_ArraySlice_l118_284_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_284 = _zz_when_ArraySlice_l118_284_1[5:0];
  assign _zz_when_ArraySlice_l173_284_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_284_1 = {1'd0, _zz_when_ArraySlice_l173_284_2};
  assign _zz_when_ArraySlice_l173_284_3 = (_zz_when_ArraySlice_l173_284_4 + _zz_when_ArraySlice_l173_284_8);
  assign _zz_when_ArraySlice_l173_284_4 = (_zz_when_ArraySlice_l173_284 - _zz_when_ArraySlice_l173_284_5);
  assign _zz_when_ArraySlice_l173_284_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_284_7);
  assign _zz_when_ArraySlice_l173_284_5 = {1'd0, _zz_when_ArraySlice_l173_284_6};
  assign _zz_when_ArraySlice_l173_284_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_284_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_285 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_285_1);
  assign _zz_when_ArraySlice_l165_285_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_285_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_285 = {1'd0, _zz_when_ArraySlice_l166_285_1};
  assign _zz_when_ArraySlice_l166_285_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_285_3);
  assign _zz_when_ArraySlice_l166_285_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_285_4);
  assign _zz_when_ArraySlice_l166_285_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_285 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_285 = (_zz_when_ArraySlice_l113_285_1 - _zz_when_ArraySlice_l113_285_4);
  assign _zz_when_ArraySlice_l113_285_1 = (_zz_when_ArraySlice_l113_285_2 + _zz_when_ArraySlice_l113_285_3);
  assign _zz_when_ArraySlice_l113_285_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_285_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_285_4 = {1'd0, _zz_when_ArraySlice_l112_285};
  assign _zz__zz_when_ArraySlice_l173_285 = (_zz__zz_when_ArraySlice_l173_285_1 + _zz__zz_when_ArraySlice_l173_285_2);
  assign _zz__zz_when_ArraySlice_l173_285_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_285_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_285_3 = {1'd0, _zz_when_ArraySlice_l112_285};
  assign _zz_when_ArraySlice_l118_285_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_285 = _zz_when_ArraySlice_l118_285_1[5:0];
  assign _zz_when_ArraySlice_l173_285_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_285_1 = {2'd0, _zz_when_ArraySlice_l173_285_2};
  assign _zz_when_ArraySlice_l173_285_3 = (_zz_when_ArraySlice_l173_285_4 + _zz_when_ArraySlice_l173_285_8);
  assign _zz_when_ArraySlice_l173_285_4 = (_zz_when_ArraySlice_l173_285 - _zz_when_ArraySlice_l173_285_5);
  assign _zz_when_ArraySlice_l173_285_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_285_7);
  assign _zz_when_ArraySlice_l173_285_5 = {1'd0, _zz_when_ArraySlice_l173_285_6};
  assign _zz_when_ArraySlice_l173_285_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_285_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_286 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_286_1);
  assign _zz_when_ArraySlice_l165_286_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_286_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_286 = {1'd0, _zz_when_ArraySlice_l166_286_1};
  assign _zz_when_ArraySlice_l166_286_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_286_3);
  assign _zz_when_ArraySlice_l166_286_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_286_4);
  assign _zz_when_ArraySlice_l166_286_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_286 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_286 = (_zz_when_ArraySlice_l113_286_1 - _zz_when_ArraySlice_l113_286_4);
  assign _zz_when_ArraySlice_l113_286_1 = (_zz_when_ArraySlice_l113_286_2 + _zz_when_ArraySlice_l113_286_3);
  assign _zz_when_ArraySlice_l113_286_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_286_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_286_4 = {1'd0, _zz_when_ArraySlice_l112_286};
  assign _zz__zz_when_ArraySlice_l173_286 = (_zz__zz_when_ArraySlice_l173_286_1 + _zz__zz_when_ArraySlice_l173_286_2);
  assign _zz__zz_when_ArraySlice_l173_286_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_286_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_286_3 = {1'd0, _zz_when_ArraySlice_l112_286};
  assign _zz_when_ArraySlice_l118_286_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_286 = _zz_when_ArraySlice_l118_286_1[5:0];
  assign _zz_when_ArraySlice_l173_286_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_286_1 = {2'd0, _zz_when_ArraySlice_l173_286_2};
  assign _zz_when_ArraySlice_l173_286_3 = (_zz_when_ArraySlice_l173_286_4 + _zz_when_ArraySlice_l173_286_8);
  assign _zz_when_ArraySlice_l173_286_4 = (_zz_when_ArraySlice_l173_286 - _zz_when_ArraySlice_l173_286_5);
  assign _zz_when_ArraySlice_l173_286_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_286_7);
  assign _zz_when_ArraySlice_l173_286_5 = {1'd0, _zz_when_ArraySlice_l173_286_6};
  assign _zz_when_ArraySlice_l173_286_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_286_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_287 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_287_1);
  assign _zz_when_ArraySlice_l165_287_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_287_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_287 = {2'd0, _zz_when_ArraySlice_l166_287_1};
  assign _zz_when_ArraySlice_l166_287_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_287_3);
  assign _zz_when_ArraySlice_l166_287_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_287_4);
  assign _zz_when_ArraySlice_l166_287_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_287 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_287 = (_zz_when_ArraySlice_l113_287_1 - _zz_when_ArraySlice_l113_287_4);
  assign _zz_when_ArraySlice_l113_287_1 = (_zz_when_ArraySlice_l113_287_2 + _zz_when_ArraySlice_l113_287_3);
  assign _zz_when_ArraySlice_l113_287_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_287_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_287_4 = {1'd0, _zz_when_ArraySlice_l112_287};
  assign _zz__zz_when_ArraySlice_l173_287 = (_zz__zz_when_ArraySlice_l173_287_1 + _zz__zz_when_ArraySlice_l173_287_2);
  assign _zz__zz_when_ArraySlice_l173_287_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_287_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_287_3 = {1'd0, _zz_when_ArraySlice_l112_287};
  assign _zz_when_ArraySlice_l118_287_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_287 = _zz_when_ArraySlice_l118_287_1[5:0];
  assign _zz_when_ArraySlice_l173_287_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_287_1 = {3'd0, _zz_when_ArraySlice_l173_287_2};
  assign _zz_when_ArraySlice_l173_287_3 = (_zz_when_ArraySlice_l173_287_4 + _zz_when_ArraySlice_l173_287_8);
  assign _zz_when_ArraySlice_l173_287_4 = (_zz_when_ArraySlice_l173_287 - _zz_when_ArraySlice_l173_287_5);
  assign _zz_when_ArraySlice_l173_287_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_287_7);
  assign _zz_when_ArraySlice_l173_287_5 = {1'd0, _zz_when_ArraySlice_l173_287_6};
  assign _zz_when_ArraySlice_l173_287_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_287_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l268_3_1 = (_zz_when_ArraySlice_l268_3_2 + _zz_when_ArraySlice_l268_3_7);
  assign _zz_when_ArraySlice_l268_3_2 = (_zz_when_ArraySlice_l268_3_3 + _zz_when_ArraySlice_l268_3_5);
  assign _zz_when_ArraySlice_l268_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l268_3_4);
  assign _zz_when_ArraySlice_l268_3_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l268_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l268_3_5 = {5'd0, _zz_when_ArraySlice_l268_3_6};
  assign _zz_when_ArraySlice_l268_3_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l268_3_7 = {1'd0, _zz_when_ArraySlice_l268_3_8};
  assign _zz_selectReadFifo_3_47 = 1'b1;
  assign _zz_selectReadFifo_3_46 = {5'd0, _zz_selectReadFifo_3_47};
  assign _zz_when_ArraySlice_l272_3_1 = (_zz_when_ArraySlice_l272_3_2 % aReg);
  assign _zz_when_ArraySlice_l272_3_2 = (handshakeTimes_3_value + _zz_when_ArraySlice_l272_3_3);
  assign _zz_when_ArraySlice_l272_3_4 = 1'b1;
  assign _zz_when_ArraySlice_l272_3_3 = {12'd0, _zz_when_ArraySlice_l272_3_4};
  assign _zz_when_ArraySlice_l276_3_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l276_3_3);
  assign _zz_when_ArraySlice_l276_3_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l276_3_3 = {1'd0, _zz_when_ArraySlice_l276_3_4};
  assign _zz_when_ArraySlice_l277_3_2 = (_zz_when_ArraySlice_l277_3_3 - _zz_when_ArraySlice_l277_3_4);
  assign _zz_when_ArraySlice_l277_3_1 = {7'd0, _zz_when_ArraySlice_l277_3_2};
  assign _zz_when_ArraySlice_l277_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l277_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l277_3_4 = {5'd0, _zz_when_ArraySlice_l277_3_5};
  assign _zz__zz_when_ArraySlice_l94_34 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_34 = (_zz_when_ArraySlice_l95_34_1 - _zz_when_ArraySlice_l95_34_4);
  assign _zz_when_ArraySlice_l95_34_1 = (_zz_when_ArraySlice_l95_34_2 + _zz_when_ArraySlice_l95_34_3);
  assign _zz_when_ArraySlice_l95_34_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_34_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_34_4 = {1'd0, _zz_when_ArraySlice_l94_34};
  assign _zz__zz_when_ArraySlice_l279_3_1 = (_zz__zz_when_ArraySlice_l279_3_2 + _zz__zz_when_ArraySlice_l279_3_3);
  assign _zz__zz_when_ArraySlice_l279_3_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l279_3_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l279_3_4 = {1'd0, _zz_when_ArraySlice_l94_34};
  assign _zz_when_ArraySlice_l99_34_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_34 = _zz_when_ArraySlice_l99_34_1[5:0];
  assign _zz_when_ArraySlice_l279_3_1 = (outSliceNumb_3_value + _zz_when_ArraySlice_l279_3_2);
  assign _zz_when_ArraySlice_l279_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l279_3_2 = {6'd0, _zz_when_ArraySlice_l279_3_3};
  assign _zz_when_ArraySlice_l279_3_4 = (_zz_when_ArraySlice_l279_3 / aReg);
  assign _zz_selectReadFifo_3_48 = (selectReadFifo_3 - _zz_selectReadFifo_3_49);
  assign _zz_selectReadFifo_3_49 = {3'd0, bReg};
  assign _zz_selectReadFifo_3_51 = 1'b1;
  assign _zz_selectReadFifo_3_50 = {5'd0, _zz_selectReadFifo_3_51};
  assign _zz_selectReadFifo_3_52 = (selectReadFifo_3 + _zz_selectReadFifo_3_53);
  assign _zz_selectReadFifo_3_53 = (3'b111 * bReg);
  assign _zz_selectReadFifo_3_55 = 1'b1;
  assign _zz_selectReadFifo_3_54 = {5'd0, _zz_selectReadFifo_3_55};
  assign _zz_when_ArraySlice_l165_288 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_288_1);
  assign _zz_when_ArraySlice_l165_288_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_288_1 = {3'd0, _zz_when_ArraySlice_l165_288_2};
  assign _zz_when_ArraySlice_l166_288 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_288_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_288_3);
  assign _zz_when_ArraySlice_l166_288_1 = {1'd0, _zz_when_ArraySlice_l166_288_2};
  assign _zz_when_ArraySlice_l166_288_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_288_4);
  assign _zz_when_ArraySlice_l166_288_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_288_4 = {3'd0, _zz_when_ArraySlice_l166_288_5};
  assign _zz__zz_when_ArraySlice_l112_288 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_288 = (_zz_when_ArraySlice_l113_288_1 - _zz_when_ArraySlice_l113_288_4);
  assign _zz_when_ArraySlice_l113_288_1 = (_zz_when_ArraySlice_l113_288_2 + _zz_when_ArraySlice_l113_288_3);
  assign _zz_when_ArraySlice_l113_288_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_288_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_288_4 = {1'd0, _zz_when_ArraySlice_l112_288};
  assign _zz__zz_when_ArraySlice_l173_288 = (_zz__zz_when_ArraySlice_l173_288_1 + _zz__zz_when_ArraySlice_l173_288_2);
  assign _zz__zz_when_ArraySlice_l173_288_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_288_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_288_3 = {1'd0, _zz_when_ArraySlice_l112_288};
  assign _zz_when_ArraySlice_l118_288_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_288 = _zz_when_ArraySlice_l118_288_1[5:0];
  assign _zz_when_ArraySlice_l173_288_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_288_2 = (_zz_when_ArraySlice_l173_288_3 + _zz_when_ArraySlice_l173_288_8);
  assign _zz_when_ArraySlice_l173_288_3 = (_zz_when_ArraySlice_l173_288 - _zz_when_ArraySlice_l173_288_4);
  assign _zz_when_ArraySlice_l173_288_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_288_6);
  assign _zz_when_ArraySlice_l173_288_4 = {1'd0, _zz_when_ArraySlice_l173_288_5};
  assign _zz_when_ArraySlice_l173_288_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_288_6 = {3'd0, _zz_when_ArraySlice_l173_288_7};
  assign _zz_when_ArraySlice_l173_288_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_289 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_289_1);
  assign _zz_when_ArraySlice_l165_289_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_289_1 = {2'd0, _zz_when_ArraySlice_l165_289_2};
  assign _zz_when_ArraySlice_l166_289 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_289_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_289_2);
  assign _zz_when_ArraySlice_l166_289_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_289_3);
  assign _zz_when_ArraySlice_l166_289_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_289_3 = {2'd0, _zz_when_ArraySlice_l166_289_4};
  assign _zz__zz_when_ArraySlice_l112_289 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_289 = (_zz_when_ArraySlice_l113_289_1 - _zz_when_ArraySlice_l113_289_4);
  assign _zz_when_ArraySlice_l113_289_1 = (_zz_when_ArraySlice_l113_289_2 + _zz_when_ArraySlice_l113_289_3);
  assign _zz_when_ArraySlice_l113_289_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_289_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_289_4 = {1'd0, _zz_when_ArraySlice_l112_289};
  assign _zz__zz_when_ArraySlice_l173_289 = (_zz__zz_when_ArraySlice_l173_289_1 + _zz__zz_when_ArraySlice_l173_289_2);
  assign _zz__zz_when_ArraySlice_l173_289_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_289_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_289_3 = {1'd0, _zz_when_ArraySlice_l112_289};
  assign _zz_when_ArraySlice_l118_289_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_289 = _zz_when_ArraySlice_l118_289_1[5:0];
  assign _zz_when_ArraySlice_l173_289_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_289_1 = {1'd0, _zz_when_ArraySlice_l173_289_2};
  assign _zz_when_ArraySlice_l173_289_3 = (_zz_when_ArraySlice_l173_289_4 + _zz_when_ArraySlice_l173_289_9);
  assign _zz_when_ArraySlice_l173_289_4 = (_zz_when_ArraySlice_l173_289 - _zz_when_ArraySlice_l173_289_5);
  assign _zz_when_ArraySlice_l173_289_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_289_7);
  assign _zz_when_ArraySlice_l173_289_5 = {1'd0, _zz_when_ArraySlice_l173_289_6};
  assign _zz_when_ArraySlice_l173_289_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_289_7 = {2'd0, _zz_when_ArraySlice_l173_289_8};
  assign _zz_when_ArraySlice_l173_289_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_290 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_290_1);
  assign _zz_when_ArraySlice_l165_290_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_290_1 = {1'd0, _zz_when_ArraySlice_l165_290_2};
  assign _zz_when_ArraySlice_l166_290 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_290_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_290_2);
  assign _zz_when_ArraySlice_l166_290_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_290_3);
  assign _zz_when_ArraySlice_l166_290_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_290_3 = {1'd0, _zz_when_ArraySlice_l166_290_4};
  assign _zz__zz_when_ArraySlice_l112_290 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_290 = (_zz_when_ArraySlice_l113_290_1 - _zz_when_ArraySlice_l113_290_4);
  assign _zz_when_ArraySlice_l113_290_1 = (_zz_when_ArraySlice_l113_290_2 + _zz_when_ArraySlice_l113_290_3);
  assign _zz_when_ArraySlice_l113_290_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_290_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_290_4 = {1'd0, _zz_when_ArraySlice_l112_290};
  assign _zz__zz_when_ArraySlice_l173_290 = (_zz__zz_when_ArraySlice_l173_290_1 + _zz__zz_when_ArraySlice_l173_290_2);
  assign _zz__zz_when_ArraySlice_l173_290_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_290_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_290_3 = {1'd0, _zz_when_ArraySlice_l112_290};
  assign _zz_when_ArraySlice_l118_290_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_290 = _zz_when_ArraySlice_l118_290_1[5:0];
  assign _zz_when_ArraySlice_l173_290_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_290_1 = {1'd0, _zz_when_ArraySlice_l173_290_2};
  assign _zz_when_ArraySlice_l173_290_3 = (_zz_when_ArraySlice_l173_290_4 + _zz_when_ArraySlice_l173_290_9);
  assign _zz_when_ArraySlice_l173_290_4 = (_zz_when_ArraySlice_l173_290 - _zz_when_ArraySlice_l173_290_5);
  assign _zz_when_ArraySlice_l173_290_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_290_7);
  assign _zz_when_ArraySlice_l173_290_5 = {1'd0, _zz_when_ArraySlice_l173_290_6};
  assign _zz_when_ArraySlice_l173_290_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_290_7 = {1'd0, _zz_when_ArraySlice_l173_290_8};
  assign _zz_when_ArraySlice_l173_290_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_291 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_291_1);
  assign _zz_when_ArraySlice_l165_291_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_291_1 = {1'd0, _zz_when_ArraySlice_l165_291_2};
  assign _zz_when_ArraySlice_l166_291 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_291_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_291_2);
  assign _zz_when_ArraySlice_l166_291_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_291_3);
  assign _zz_when_ArraySlice_l166_291_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_291_3 = {1'd0, _zz_when_ArraySlice_l166_291_4};
  assign _zz__zz_when_ArraySlice_l112_291 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_291 = (_zz_when_ArraySlice_l113_291_1 - _zz_when_ArraySlice_l113_291_4);
  assign _zz_when_ArraySlice_l113_291_1 = (_zz_when_ArraySlice_l113_291_2 + _zz_when_ArraySlice_l113_291_3);
  assign _zz_when_ArraySlice_l113_291_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_291_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_291_4 = {1'd0, _zz_when_ArraySlice_l112_291};
  assign _zz__zz_when_ArraySlice_l173_291 = (_zz__zz_when_ArraySlice_l173_291_1 + _zz__zz_when_ArraySlice_l173_291_2);
  assign _zz__zz_when_ArraySlice_l173_291_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_291_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_291_3 = {1'd0, _zz_when_ArraySlice_l112_291};
  assign _zz_when_ArraySlice_l118_291_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_291 = _zz_when_ArraySlice_l118_291_1[5:0];
  assign _zz_when_ArraySlice_l173_291_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_291_1 = {1'd0, _zz_when_ArraySlice_l173_291_2};
  assign _zz_when_ArraySlice_l173_291_3 = (_zz_when_ArraySlice_l173_291_4 + _zz_when_ArraySlice_l173_291_9);
  assign _zz_when_ArraySlice_l173_291_4 = (_zz_when_ArraySlice_l173_291 - _zz_when_ArraySlice_l173_291_5);
  assign _zz_when_ArraySlice_l173_291_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_291_7);
  assign _zz_when_ArraySlice_l173_291_5 = {1'd0, _zz_when_ArraySlice_l173_291_6};
  assign _zz_when_ArraySlice_l173_291_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_291_7 = {1'd0, _zz_when_ArraySlice_l173_291_8};
  assign _zz_when_ArraySlice_l173_291_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_292 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_292_1);
  assign _zz_when_ArraySlice_l165_292_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_292 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_292_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_292_2);
  assign _zz_when_ArraySlice_l166_292_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_292_3);
  assign _zz_when_ArraySlice_l166_292_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_292 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_292 = (_zz_when_ArraySlice_l113_292_1 - _zz_when_ArraySlice_l113_292_4);
  assign _zz_when_ArraySlice_l113_292_1 = (_zz_when_ArraySlice_l113_292_2 + _zz_when_ArraySlice_l113_292_3);
  assign _zz_when_ArraySlice_l113_292_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_292_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_292_4 = {1'd0, _zz_when_ArraySlice_l112_292};
  assign _zz__zz_when_ArraySlice_l173_292 = (_zz__zz_when_ArraySlice_l173_292_1 + _zz__zz_when_ArraySlice_l173_292_2);
  assign _zz__zz_when_ArraySlice_l173_292_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_292_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_292_3 = {1'd0, _zz_when_ArraySlice_l112_292};
  assign _zz_when_ArraySlice_l118_292_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_292 = _zz_when_ArraySlice_l118_292_1[5:0];
  assign _zz_when_ArraySlice_l173_292_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_292_1 = {1'd0, _zz_when_ArraySlice_l173_292_2};
  assign _zz_when_ArraySlice_l173_292_3 = (_zz_when_ArraySlice_l173_292_4 + _zz_when_ArraySlice_l173_292_8);
  assign _zz_when_ArraySlice_l173_292_4 = (_zz_when_ArraySlice_l173_292 - _zz_when_ArraySlice_l173_292_5);
  assign _zz_when_ArraySlice_l173_292_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_292_7);
  assign _zz_when_ArraySlice_l173_292_5 = {1'd0, _zz_when_ArraySlice_l173_292_6};
  assign _zz_when_ArraySlice_l173_292_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_292_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_293 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_293_1);
  assign _zz_when_ArraySlice_l165_293_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_293_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_293 = {1'd0, _zz_when_ArraySlice_l166_293_1};
  assign _zz_when_ArraySlice_l166_293_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_293_3);
  assign _zz_when_ArraySlice_l166_293_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_293_4);
  assign _zz_when_ArraySlice_l166_293_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_293 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_293 = (_zz_when_ArraySlice_l113_293_1 - _zz_when_ArraySlice_l113_293_4);
  assign _zz_when_ArraySlice_l113_293_1 = (_zz_when_ArraySlice_l113_293_2 + _zz_when_ArraySlice_l113_293_3);
  assign _zz_when_ArraySlice_l113_293_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_293_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_293_4 = {1'd0, _zz_when_ArraySlice_l112_293};
  assign _zz__zz_when_ArraySlice_l173_293 = (_zz__zz_when_ArraySlice_l173_293_1 + _zz__zz_when_ArraySlice_l173_293_2);
  assign _zz__zz_when_ArraySlice_l173_293_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_293_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_293_3 = {1'd0, _zz_when_ArraySlice_l112_293};
  assign _zz_when_ArraySlice_l118_293_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_293 = _zz_when_ArraySlice_l118_293_1[5:0];
  assign _zz_when_ArraySlice_l173_293_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_293_1 = {2'd0, _zz_when_ArraySlice_l173_293_2};
  assign _zz_when_ArraySlice_l173_293_3 = (_zz_when_ArraySlice_l173_293_4 + _zz_when_ArraySlice_l173_293_8);
  assign _zz_when_ArraySlice_l173_293_4 = (_zz_when_ArraySlice_l173_293 - _zz_when_ArraySlice_l173_293_5);
  assign _zz_when_ArraySlice_l173_293_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_293_7);
  assign _zz_when_ArraySlice_l173_293_5 = {1'd0, _zz_when_ArraySlice_l173_293_6};
  assign _zz_when_ArraySlice_l173_293_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_293_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_294 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_294_1);
  assign _zz_when_ArraySlice_l165_294_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_294_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_294 = {1'd0, _zz_when_ArraySlice_l166_294_1};
  assign _zz_when_ArraySlice_l166_294_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_294_3);
  assign _zz_when_ArraySlice_l166_294_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_294_4);
  assign _zz_when_ArraySlice_l166_294_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_294 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_294 = (_zz_when_ArraySlice_l113_294_1 - _zz_when_ArraySlice_l113_294_4);
  assign _zz_when_ArraySlice_l113_294_1 = (_zz_when_ArraySlice_l113_294_2 + _zz_when_ArraySlice_l113_294_3);
  assign _zz_when_ArraySlice_l113_294_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_294_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_294_4 = {1'd0, _zz_when_ArraySlice_l112_294};
  assign _zz__zz_when_ArraySlice_l173_294 = (_zz__zz_when_ArraySlice_l173_294_1 + _zz__zz_when_ArraySlice_l173_294_2);
  assign _zz__zz_when_ArraySlice_l173_294_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_294_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_294_3 = {1'd0, _zz_when_ArraySlice_l112_294};
  assign _zz_when_ArraySlice_l118_294_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_294 = _zz_when_ArraySlice_l118_294_1[5:0];
  assign _zz_when_ArraySlice_l173_294_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_294_1 = {2'd0, _zz_when_ArraySlice_l173_294_2};
  assign _zz_when_ArraySlice_l173_294_3 = (_zz_when_ArraySlice_l173_294_4 + _zz_when_ArraySlice_l173_294_8);
  assign _zz_when_ArraySlice_l173_294_4 = (_zz_when_ArraySlice_l173_294 - _zz_when_ArraySlice_l173_294_5);
  assign _zz_when_ArraySlice_l173_294_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_294_7);
  assign _zz_when_ArraySlice_l173_294_5 = {1'd0, _zz_when_ArraySlice_l173_294_6};
  assign _zz_when_ArraySlice_l173_294_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_294_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_295 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_295_1);
  assign _zz_when_ArraySlice_l165_295_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_295_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_295 = {2'd0, _zz_when_ArraySlice_l166_295_1};
  assign _zz_when_ArraySlice_l166_295_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_295_3);
  assign _zz_when_ArraySlice_l166_295_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_295_4);
  assign _zz_when_ArraySlice_l166_295_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_295 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_295 = (_zz_when_ArraySlice_l113_295_1 - _zz_when_ArraySlice_l113_295_4);
  assign _zz_when_ArraySlice_l113_295_1 = (_zz_when_ArraySlice_l113_295_2 + _zz_when_ArraySlice_l113_295_3);
  assign _zz_when_ArraySlice_l113_295_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_295_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_295_4 = {1'd0, _zz_when_ArraySlice_l112_295};
  assign _zz__zz_when_ArraySlice_l173_295 = (_zz__zz_when_ArraySlice_l173_295_1 + _zz__zz_when_ArraySlice_l173_295_2);
  assign _zz__zz_when_ArraySlice_l173_295_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_295_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_295_3 = {1'd0, _zz_when_ArraySlice_l112_295};
  assign _zz_when_ArraySlice_l118_295_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_295 = _zz_when_ArraySlice_l118_295_1[5:0];
  assign _zz_when_ArraySlice_l173_295_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_295_1 = {3'd0, _zz_when_ArraySlice_l173_295_2};
  assign _zz_when_ArraySlice_l173_295_3 = (_zz_when_ArraySlice_l173_295_4 + _zz_when_ArraySlice_l173_295_8);
  assign _zz_when_ArraySlice_l173_295_4 = (_zz_when_ArraySlice_l173_295 - _zz_when_ArraySlice_l173_295_5);
  assign _zz_when_ArraySlice_l173_295_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_295_7);
  assign _zz_when_ArraySlice_l173_295_5 = {1'd0, _zz_when_ArraySlice_l173_295_6};
  assign _zz_when_ArraySlice_l173_295_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_295_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l288_3_1 = (_zz_when_ArraySlice_l288_3_2 + _zz_when_ArraySlice_l288_3_7);
  assign _zz_when_ArraySlice_l288_3_2 = (_zz_when_ArraySlice_l288_3_3 + _zz_when_ArraySlice_l288_3_5);
  assign _zz_when_ArraySlice_l288_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l288_3_4);
  assign _zz_when_ArraySlice_l288_3_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l288_3_5 = {5'd0, _zz_when_ArraySlice_l288_3_6};
  assign _zz_when_ArraySlice_l288_3_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l288_3_7 = {1'd0, _zz_when_ArraySlice_l288_3_8};
  assign _zz_selectReadFifo_3_57 = 1'b1;
  assign _zz_selectReadFifo_3_56 = {5'd0, _zz_selectReadFifo_3_57};
  assign _zz_when_ArraySlice_l292_3_1 = (_zz_when_ArraySlice_l292_3_2 % aReg);
  assign _zz_when_ArraySlice_l292_3_2 = (handshakeTimes_3_value + _zz_when_ArraySlice_l292_3_3);
  assign _zz_when_ArraySlice_l292_3_4 = 1'b1;
  assign _zz_when_ArraySlice_l292_3_3 = {12'd0, _zz_when_ArraySlice_l292_3_4};
  assign _zz_when_ArraySlice_l303_3_2 = (_zz_when_ArraySlice_l303_3_3 - _zz_when_ArraySlice_l303_3_4);
  assign _zz_when_ArraySlice_l303_3_1 = {7'd0, _zz_when_ArraySlice_l303_3_2};
  assign _zz_when_ArraySlice_l303_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l303_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l303_3_4 = {5'd0, _zz_when_ArraySlice_l303_3_5};
  assign _zz__zz_when_ArraySlice_l94_35 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_35 = (_zz_when_ArraySlice_l95_35_1 - _zz_when_ArraySlice_l95_35_4);
  assign _zz_when_ArraySlice_l95_35_1 = (_zz_when_ArraySlice_l95_35_2 + _zz_when_ArraySlice_l95_35_3);
  assign _zz_when_ArraySlice_l95_35_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_35_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_35_4 = {1'd0, _zz_when_ArraySlice_l94_35};
  assign _zz__zz_when_ArraySlice_l304_3_1 = (_zz__zz_when_ArraySlice_l304_3_2 + _zz__zz_when_ArraySlice_l304_3_3);
  assign _zz__zz_when_ArraySlice_l304_3_2 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l304_3_3 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l304_3_4 = {1'd0, _zz_when_ArraySlice_l94_35};
  assign _zz_when_ArraySlice_l99_35_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_35 = _zz_when_ArraySlice_l99_35_1[5:0];
  assign _zz_when_ArraySlice_l304_3_1 = (outSliceNumb_3_value + _zz_when_ArraySlice_l304_3_2);
  assign _zz_when_ArraySlice_l304_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l304_3_2 = {6'd0, _zz_when_ArraySlice_l304_3_3};
  assign _zz_when_ArraySlice_l304_3_4 = (_zz_when_ArraySlice_l304_3 / aReg);
  assign _zz_selectReadFifo_3_58 = (selectReadFifo_3 - _zz_selectReadFifo_3_59);
  assign _zz_selectReadFifo_3_59 = {3'd0, bReg};
  assign _zz_selectReadFifo_3_61 = 1'b1;
  assign _zz_selectReadFifo_3_60 = {5'd0, _zz_selectReadFifo_3_61};
  assign _zz_when_ArraySlice_l165_296 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_296_1);
  assign _zz_when_ArraySlice_l165_296_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_296_1 = {3'd0, _zz_when_ArraySlice_l165_296_2};
  assign _zz_when_ArraySlice_l166_296 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_296_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_296_3);
  assign _zz_when_ArraySlice_l166_296_1 = {1'd0, _zz_when_ArraySlice_l166_296_2};
  assign _zz_when_ArraySlice_l166_296_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_296_4);
  assign _zz_when_ArraySlice_l166_296_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_296_4 = {3'd0, _zz_when_ArraySlice_l166_296_5};
  assign _zz__zz_when_ArraySlice_l112_296 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_296 = (_zz_when_ArraySlice_l113_296_1 - _zz_when_ArraySlice_l113_296_4);
  assign _zz_when_ArraySlice_l113_296_1 = (_zz_when_ArraySlice_l113_296_2 + _zz_when_ArraySlice_l113_296_3);
  assign _zz_when_ArraySlice_l113_296_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_296_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_296_4 = {1'd0, _zz_when_ArraySlice_l112_296};
  assign _zz__zz_when_ArraySlice_l173_296 = (_zz__zz_when_ArraySlice_l173_296_1 + _zz__zz_when_ArraySlice_l173_296_2);
  assign _zz__zz_when_ArraySlice_l173_296_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_296_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_296_3 = {1'd0, _zz_when_ArraySlice_l112_296};
  assign _zz_when_ArraySlice_l118_296_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_296 = _zz_when_ArraySlice_l118_296_1[5:0];
  assign _zz_when_ArraySlice_l173_296_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_296_2 = (_zz_when_ArraySlice_l173_296_3 + _zz_when_ArraySlice_l173_296_8);
  assign _zz_when_ArraySlice_l173_296_3 = (_zz_when_ArraySlice_l173_296 - _zz_when_ArraySlice_l173_296_4);
  assign _zz_when_ArraySlice_l173_296_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_296_6);
  assign _zz_when_ArraySlice_l173_296_4 = {1'd0, _zz_when_ArraySlice_l173_296_5};
  assign _zz_when_ArraySlice_l173_296_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_296_6 = {3'd0, _zz_when_ArraySlice_l173_296_7};
  assign _zz_when_ArraySlice_l173_296_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_297 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_297_1);
  assign _zz_when_ArraySlice_l165_297_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_297_1 = {2'd0, _zz_when_ArraySlice_l165_297_2};
  assign _zz_when_ArraySlice_l166_297 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_297_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_297_2);
  assign _zz_when_ArraySlice_l166_297_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_297_3);
  assign _zz_when_ArraySlice_l166_297_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_297_3 = {2'd0, _zz_when_ArraySlice_l166_297_4};
  assign _zz__zz_when_ArraySlice_l112_297 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_297 = (_zz_when_ArraySlice_l113_297_1 - _zz_when_ArraySlice_l113_297_4);
  assign _zz_when_ArraySlice_l113_297_1 = (_zz_when_ArraySlice_l113_297_2 + _zz_when_ArraySlice_l113_297_3);
  assign _zz_when_ArraySlice_l113_297_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_297_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_297_4 = {1'd0, _zz_when_ArraySlice_l112_297};
  assign _zz__zz_when_ArraySlice_l173_297 = (_zz__zz_when_ArraySlice_l173_297_1 + _zz__zz_when_ArraySlice_l173_297_2);
  assign _zz__zz_when_ArraySlice_l173_297_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_297_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_297_3 = {1'd0, _zz_when_ArraySlice_l112_297};
  assign _zz_when_ArraySlice_l118_297_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_297 = _zz_when_ArraySlice_l118_297_1[5:0];
  assign _zz_when_ArraySlice_l173_297_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_297_1 = {1'd0, _zz_when_ArraySlice_l173_297_2};
  assign _zz_when_ArraySlice_l173_297_3 = (_zz_when_ArraySlice_l173_297_4 + _zz_when_ArraySlice_l173_297_9);
  assign _zz_when_ArraySlice_l173_297_4 = (_zz_when_ArraySlice_l173_297 - _zz_when_ArraySlice_l173_297_5);
  assign _zz_when_ArraySlice_l173_297_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_297_7);
  assign _zz_when_ArraySlice_l173_297_5 = {1'd0, _zz_when_ArraySlice_l173_297_6};
  assign _zz_when_ArraySlice_l173_297_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_297_7 = {2'd0, _zz_when_ArraySlice_l173_297_8};
  assign _zz_when_ArraySlice_l173_297_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_298 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_298_1);
  assign _zz_when_ArraySlice_l165_298_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_298_1 = {1'd0, _zz_when_ArraySlice_l165_298_2};
  assign _zz_when_ArraySlice_l166_298 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_298_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_298_2);
  assign _zz_when_ArraySlice_l166_298_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_298_3);
  assign _zz_when_ArraySlice_l166_298_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_298_3 = {1'd0, _zz_when_ArraySlice_l166_298_4};
  assign _zz__zz_when_ArraySlice_l112_298 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_298 = (_zz_when_ArraySlice_l113_298_1 - _zz_when_ArraySlice_l113_298_4);
  assign _zz_when_ArraySlice_l113_298_1 = (_zz_when_ArraySlice_l113_298_2 + _zz_when_ArraySlice_l113_298_3);
  assign _zz_when_ArraySlice_l113_298_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_298_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_298_4 = {1'd0, _zz_when_ArraySlice_l112_298};
  assign _zz__zz_when_ArraySlice_l173_298 = (_zz__zz_when_ArraySlice_l173_298_1 + _zz__zz_when_ArraySlice_l173_298_2);
  assign _zz__zz_when_ArraySlice_l173_298_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_298_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_298_3 = {1'd0, _zz_when_ArraySlice_l112_298};
  assign _zz_when_ArraySlice_l118_298_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_298 = _zz_when_ArraySlice_l118_298_1[5:0];
  assign _zz_when_ArraySlice_l173_298_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_298_1 = {1'd0, _zz_when_ArraySlice_l173_298_2};
  assign _zz_when_ArraySlice_l173_298_3 = (_zz_when_ArraySlice_l173_298_4 + _zz_when_ArraySlice_l173_298_9);
  assign _zz_when_ArraySlice_l173_298_4 = (_zz_when_ArraySlice_l173_298 - _zz_when_ArraySlice_l173_298_5);
  assign _zz_when_ArraySlice_l173_298_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_298_7);
  assign _zz_when_ArraySlice_l173_298_5 = {1'd0, _zz_when_ArraySlice_l173_298_6};
  assign _zz_when_ArraySlice_l173_298_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_298_7 = {1'd0, _zz_when_ArraySlice_l173_298_8};
  assign _zz_when_ArraySlice_l173_298_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_299 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_299_1);
  assign _zz_when_ArraySlice_l165_299_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_299_1 = {1'd0, _zz_when_ArraySlice_l165_299_2};
  assign _zz_when_ArraySlice_l166_299 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_299_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_299_2);
  assign _zz_when_ArraySlice_l166_299_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_299_3);
  assign _zz_when_ArraySlice_l166_299_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_299_3 = {1'd0, _zz_when_ArraySlice_l166_299_4};
  assign _zz__zz_when_ArraySlice_l112_299 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_299 = (_zz_when_ArraySlice_l113_299_1 - _zz_when_ArraySlice_l113_299_4);
  assign _zz_when_ArraySlice_l113_299_1 = (_zz_when_ArraySlice_l113_299_2 + _zz_when_ArraySlice_l113_299_3);
  assign _zz_when_ArraySlice_l113_299_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_299_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_299_4 = {1'd0, _zz_when_ArraySlice_l112_299};
  assign _zz__zz_when_ArraySlice_l173_299 = (_zz__zz_when_ArraySlice_l173_299_1 + _zz__zz_when_ArraySlice_l173_299_2);
  assign _zz__zz_when_ArraySlice_l173_299_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_299_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_299_3 = {1'd0, _zz_when_ArraySlice_l112_299};
  assign _zz_when_ArraySlice_l118_299_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_299 = _zz_when_ArraySlice_l118_299_1[5:0];
  assign _zz_when_ArraySlice_l173_299_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_299_1 = {1'd0, _zz_when_ArraySlice_l173_299_2};
  assign _zz_when_ArraySlice_l173_299_3 = (_zz_when_ArraySlice_l173_299_4 + _zz_when_ArraySlice_l173_299_9);
  assign _zz_when_ArraySlice_l173_299_4 = (_zz_when_ArraySlice_l173_299 - _zz_when_ArraySlice_l173_299_5);
  assign _zz_when_ArraySlice_l173_299_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_299_7);
  assign _zz_when_ArraySlice_l173_299_5 = {1'd0, _zz_when_ArraySlice_l173_299_6};
  assign _zz_when_ArraySlice_l173_299_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_299_7 = {1'd0, _zz_when_ArraySlice_l173_299_8};
  assign _zz_when_ArraySlice_l173_299_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_300 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_300_1);
  assign _zz_when_ArraySlice_l165_300_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_300 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_300_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_300_2);
  assign _zz_when_ArraySlice_l166_300_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_300_3);
  assign _zz_when_ArraySlice_l166_300_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_300 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_300 = (_zz_when_ArraySlice_l113_300_1 - _zz_when_ArraySlice_l113_300_4);
  assign _zz_when_ArraySlice_l113_300_1 = (_zz_when_ArraySlice_l113_300_2 + _zz_when_ArraySlice_l113_300_3);
  assign _zz_when_ArraySlice_l113_300_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_300_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_300_4 = {1'd0, _zz_when_ArraySlice_l112_300};
  assign _zz__zz_when_ArraySlice_l173_300 = (_zz__zz_when_ArraySlice_l173_300_1 + _zz__zz_when_ArraySlice_l173_300_2);
  assign _zz__zz_when_ArraySlice_l173_300_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_300_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_300_3 = {1'd0, _zz_when_ArraySlice_l112_300};
  assign _zz_when_ArraySlice_l118_300_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_300 = _zz_when_ArraySlice_l118_300_1[5:0];
  assign _zz_when_ArraySlice_l173_300_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_300_1 = {1'd0, _zz_when_ArraySlice_l173_300_2};
  assign _zz_when_ArraySlice_l173_300_3 = (_zz_when_ArraySlice_l173_300_4 + _zz_when_ArraySlice_l173_300_8);
  assign _zz_when_ArraySlice_l173_300_4 = (_zz_when_ArraySlice_l173_300 - _zz_when_ArraySlice_l173_300_5);
  assign _zz_when_ArraySlice_l173_300_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_300_7);
  assign _zz_when_ArraySlice_l173_300_5 = {1'd0, _zz_when_ArraySlice_l173_300_6};
  assign _zz_when_ArraySlice_l173_300_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_300_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_301 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_301_1);
  assign _zz_when_ArraySlice_l165_301_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_301_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_301 = {1'd0, _zz_when_ArraySlice_l166_301_1};
  assign _zz_when_ArraySlice_l166_301_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_301_3);
  assign _zz_when_ArraySlice_l166_301_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_301_4);
  assign _zz_when_ArraySlice_l166_301_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_301 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_301 = (_zz_when_ArraySlice_l113_301_1 - _zz_when_ArraySlice_l113_301_4);
  assign _zz_when_ArraySlice_l113_301_1 = (_zz_when_ArraySlice_l113_301_2 + _zz_when_ArraySlice_l113_301_3);
  assign _zz_when_ArraySlice_l113_301_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_301_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_301_4 = {1'd0, _zz_when_ArraySlice_l112_301};
  assign _zz__zz_when_ArraySlice_l173_301 = (_zz__zz_when_ArraySlice_l173_301_1 + _zz__zz_when_ArraySlice_l173_301_2);
  assign _zz__zz_when_ArraySlice_l173_301_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_301_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_301_3 = {1'd0, _zz_when_ArraySlice_l112_301};
  assign _zz_when_ArraySlice_l118_301_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_301 = _zz_when_ArraySlice_l118_301_1[5:0];
  assign _zz_when_ArraySlice_l173_301_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_301_1 = {2'd0, _zz_when_ArraySlice_l173_301_2};
  assign _zz_when_ArraySlice_l173_301_3 = (_zz_when_ArraySlice_l173_301_4 + _zz_when_ArraySlice_l173_301_8);
  assign _zz_when_ArraySlice_l173_301_4 = (_zz_when_ArraySlice_l173_301 - _zz_when_ArraySlice_l173_301_5);
  assign _zz_when_ArraySlice_l173_301_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_301_7);
  assign _zz_when_ArraySlice_l173_301_5 = {1'd0, _zz_when_ArraySlice_l173_301_6};
  assign _zz_when_ArraySlice_l173_301_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_301_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_302 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_302_1);
  assign _zz_when_ArraySlice_l165_302_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_302_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_302 = {1'd0, _zz_when_ArraySlice_l166_302_1};
  assign _zz_when_ArraySlice_l166_302_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_302_3);
  assign _zz_when_ArraySlice_l166_302_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_302_4);
  assign _zz_when_ArraySlice_l166_302_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_302 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_302 = (_zz_when_ArraySlice_l113_302_1 - _zz_when_ArraySlice_l113_302_4);
  assign _zz_when_ArraySlice_l113_302_1 = (_zz_when_ArraySlice_l113_302_2 + _zz_when_ArraySlice_l113_302_3);
  assign _zz_when_ArraySlice_l113_302_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_302_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_302_4 = {1'd0, _zz_when_ArraySlice_l112_302};
  assign _zz__zz_when_ArraySlice_l173_302 = (_zz__zz_when_ArraySlice_l173_302_1 + _zz__zz_when_ArraySlice_l173_302_2);
  assign _zz__zz_when_ArraySlice_l173_302_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_302_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_302_3 = {1'd0, _zz_when_ArraySlice_l112_302};
  assign _zz_when_ArraySlice_l118_302_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_302 = _zz_when_ArraySlice_l118_302_1[5:0];
  assign _zz_when_ArraySlice_l173_302_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_302_1 = {2'd0, _zz_when_ArraySlice_l173_302_2};
  assign _zz_when_ArraySlice_l173_302_3 = (_zz_when_ArraySlice_l173_302_4 + _zz_when_ArraySlice_l173_302_8);
  assign _zz_when_ArraySlice_l173_302_4 = (_zz_when_ArraySlice_l173_302 - _zz_when_ArraySlice_l173_302_5);
  assign _zz_when_ArraySlice_l173_302_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_302_7);
  assign _zz_when_ArraySlice_l173_302_5 = {1'd0, _zz_when_ArraySlice_l173_302_6};
  assign _zz_when_ArraySlice_l173_302_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_302_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_303 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_303_1);
  assign _zz_when_ArraySlice_l165_303_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_303_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_303 = {2'd0, _zz_when_ArraySlice_l166_303_1};
  assign _zz_when_ArraySlice_l166_303_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_303_3);
  assign _zz_when_ArraySlice_l166_303_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_303_4);
  assign _zz_when_ArraySlice_l166_303_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_303 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_303 = (_zz_when_ArraySlice_l113_303_1 - _zz_when_ArraySlice_l113_303_4);
  assign _zz_when_ArraySlice_l113_303_1 = (_zz_when_ArraySlice_l113_303_2 + _zz_when_ArraySlice_l113_303_3);
  assign _zz_when_ArraySlice_l113_303_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_303_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_303_4 = {1'd0, _zz_when_ArraySlice_l112_303};
  assign _zz__zz_when_ArraySlice_l173_303 = (_zz__zz_when_ArraySlice_l173_303_1 + _zz__zz_when_ArraySlice_l173_303_2);
  assign _zz__zz_when_ArraySlice_l173_303_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_303_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_303_3 = {1'd0, _zz_when_ArraySlice_l112_303};
  assign _zz_when_ArraySlice_l118_303_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_303 = _zz_when_ArraySlice_l118_303_1[5:0];
  assign _zz_when_ArraySlice_l173_303_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_303_1 = {3'd0, _zz_when_ArraySlice_l173_303_2};
  assign _zz_when_ArraySlice_l173_303_3 = (_zz_when_ArraySlice_l173_303_4 + _zz_when_ArraySlice_l173_303_8);
  assign _zz_when_ArraySlice_l173_303_4 = (_zz_when_ArraySlice_l173_303 - _zz_when_ArraySlice_l173_303_5);
  assign _zz_when_ArraySlice_l173_303_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_303_7);
  assign _zz_when_ArraySlice_l173_303_5 = {1'd0, _zz_when_ArraySlice_l173_303_6};
  assign _zz_when_ArraySlice_l173_303_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_303_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_3_63 = 1'b1;
  assign _zz_selectReadFifo_3_62 = {5'd0, _zz_selectReadFifo_3_63};
  assign _zz_when_ArraySlice_l315_3_1 = (_zz_when_ArraySlice_l315_3_2 % aReg);
  assign _zz_when_ArraySlice_l315_3_2 = (handshakeTimes_3_value + _zz_when_ArraySlice_l315_3_3);
  assign _zz_when_ArraySlice_l315_3_4 = 1'b1;
  assign _zz_when_ArraySlice_l315_3_3 = {12'd0, _zz_when_ArraySlice_l315_3_4};
  assign _zz_when_ArraySlice_l301_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l301_3_1);
  assign _zz_when_ArraySlice_l301_3_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l301_3_1 = {1'd0, _zz_when_ArraySlice_l301_3_2};
  assign _zz_when_ArraySlice_l322_3_2 = (_zz_when_ArraySlice_l322_3_3 - _zz_when_ArraySlice_l322_3_4);
  assign _zz_when_ArraySlice_l322_3_1 = {7'd0, _zz_when_ArraySlice_l322_3_2};
  assign _zz_when_ArraySlice_l322_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l322_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l322_3_4 = {5'd0, _zz_when_ArraySlice_l322_3_5};
  assign _zz_when_ArraySlice_l240_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l240_4_1);
  assign _zz_when_ArraySlice_l240_4_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l241_4_1 = (selectReadFifo_4 + _zz_when_ArraySlice_l241_4_2);
  assign _zz_when_ArraySlice_l241_4_2 = (bReg * 3'b100);
  assign _zz__zz_outputStreamArrayData_4_valid_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l247_4_2 = 1'b1;
  assign _zz_when_ArraySlice_l247_4_1 = {6'd0, _zz_when_ArraySlice_l247_4_2};
  assign _zz_when_ArraySlice_l247_4_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l247_4_5);
  assign _zz_when_ArraySlice_l247_4_5 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l248_4_2 = (_zz_when_ArraySlice_l248_4_3 - _zz_when_ArraySlice_l248_4_4);
  assign _zz_when_ArraySlice_l248_4_1 = {7'd0, _zz_when_ArraySlice_l248_4_2};
  assign _zz_when_ArraySlice_l248_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l248_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l248_4_4 = {5'd0, _zz_when_ArraySlice_l248_4_5};
  assign _zz_selectReadFifo_4_32 = (selectReadFifo_4 - _zz_selectReadFifo_4_33);
  assign _zz_selectReadFifo_4_33 = {3'd0, bReg};
  assign _zz_selectReadFifo_4_35 = 1'b1;
  assign _zz_selectReadFifo_4_34 = {5'd0, _zz_selectReadFifo_4_35};
  assign _zz_selectReadFifo_4_37 = 1'b1;
  assign _zz_selectReadFifo_4_36 = {5'd0, _zz_selectReadFifo_4_37};
  assign _zz_when_ArraySlice_l251_4 = (_zz_when_ArraySlice_l251_4_1 % aReg);
  assign _zz_when_ArraySlice_l251_4_1 = (handshakeTimes_4_value + _zz_when_ArraySlice_l251_4_2);
  assign _zz_when_ArraySlice_l251_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l251_4_2 = {12'd0, _zz_when_ArraySlice_l251_4_3};
  assign _zz_when_ArraySlice_l256_4_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l256_4_3);
  assign _zz_when_ArraySlice_l256_4_3 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l256_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l256_4_4 = {6'd0, _zz_when_ArraySlice_l256_4_5};
  assign _zz_when_ArraySlice_l257_4_2 = (_zz_when_ArraySlice_l257_4_3 - _zz_when_ArraySlice_l257_4_4);
  assign _zz_when_ArraySlice_l257_4_1 = {7'd0, _zz_when_ArraySlice_l257_4_2};
  assign _zz_when_ArraySlice_l257_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l257_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l257_4_4 = {5'd0, _zz_when_ArraySlice_l257_4_5};
  assign _zz__zz_when_ArraySlice_l94_36 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_36 = (_zz_when_ArraySlice_l95_36_1 - _zz_when_ArraySlice_l95_36_4);
  assign _zz_when_ArraySlice_l95_36_1 = (_zz_when_ArraySlice_l95_36_2 + _zz_when_ArraySlice_l95_36_3);
  assign _zz_when_ArraySlice_l95_36_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_36_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_36_4 = {1'd0, _zz_when_ArraySlice_l94_36};
  assign _zz__zz_when_ArraySlice_l259_4 = (_zz__zz_when_ArraySlice_l259_4_1 + _zz__zz_when_ArraySlice_l259_4_2);
  assign _zz__zz_when_ArraySlice_l259_4_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l259_4_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l259_4_3 = {1'd0, _zz_when_ArraySlice_l94_36};
  assign _zz_when_ArraySlice_l99_36_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_36 = _zz_when_ArraySlice_l99_36_1[5:0];
  assign _zz_when_ArraySlice_l259_4_1 = (outSliceNumb_4_value + _zz_when_ArraySlice_l259_4_2);
  assign _zz_when_ArraySlice_l259_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l259_4_2 = {6'd0, _zz_when_ArraySlice_l259_4_3};
  assign _zz_when_ArraySlice_l259_4_4 = (_zz_when_ArraySlice_l259_4 / aReg);
  assign _zz_selectReadFifo_4_38 = (selectReadFifo_4 - _zz_selectReadFifo_4_39);
  assign _zz_selectReadFifo_4_39 = {3'd0, bReg};
  assign _zz_selectReadFifo_4_41 = 1'b1;
  assign _zz_selectReadFifo_4_40 = {5'd0, _zz_selectReadFifo_4_41};
  assign _zz_selectReadFifo_4_42 = (selectReadFifo_4 + _zz_selectReadFifo_4_43);
  assign _zz_selectReadFifo_4_43 = (3'b111 * bReg);
  assign _zz_selectReadFifo_4_45 = 1'b1;
  assign _zz_selectReadFifo_4_44 = {5'd0, _zz_selectReadFifo_4_45};
  assign _zz_when_ArraySlice_l165_304 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_304_1);
  assign _zz_when_ArraySlice_l165_304_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_304_1 = {3'd0, _zz_when_ArraySlice_l165_304_2};
  assign _zz_when_ArraySlice_l166_304 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_304_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_304_3);
  assign _zz_when_ArraySlice_l166_304_1 = {1'd0, _zz_when_ArraySlice_l166_304_2};
  assign _zz_when_ArraySlice_l166_304_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_304_4);
  assign _zz_when_ArraySlice_l166_304_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_304_4 = {3'd0, _zz_when_ArraySlice_l166_304_5};
  assign _zz__zz_when_ArraySlice_l112_304 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_304 = (_zz_when_ArraySlice_l113_304_1 - _zz_when_ArraySlice_l113_304_4);
  assign _zz_when_ArraySlice_l113_304_1 = (_zz_when_ArraySlice_l113_304_2 + _zz_when_ArraySlice_l113_304_3);
  assign _zz_when_ArraySlice_l113_304_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_304_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_304_4 = {1'd0, _zz_when_ArraySlice_l112_304};
  assign _zz__zz_when_ArraySlice_l173_304 = (_zz__zz_when_ArraySlice_l173_304_1 + _zz__zz_when_ArraySlice_l173_304_2);
  assign _zz__zz_when_ArraySlice_l173_304_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_304_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_304_3 = {1'd0, _zz_when_ArraySlice_l112_304};
  assign _zz_when_ArraySlice_l118_304_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_304 = _zz_when_ArraySlice_l118_304_1[5:0];
  assign _zz_when_ArraySlice_l173_304_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_304_2 = (_zz_when_ArraySlice_l173_304_3 + _zz_when_ArraySlice_l173_304_8);
  assign _zz_when_ArraySlice_l173_304_3 = (_zz_when_ArraySlice_l173_304 - _zz_when_ArraySlice_l173_304_4);
  assign _zz_when_ArraySlice_l173_304_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_304_6);
  assign _zz_when_ArraySlice_l173_304_4 = {1'd0, _zz_when_ArraySlice_l173_304_5};
  assign _zz_when_ArraySlice_l173_304_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_304_6 = {3'd0, _zz_when_ArraySlice_l173_304_7};
  assign _zz_when_ArraySlice_l173_304_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_305 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_305_1);
  assign _zz_when_ArraySlice_l165_305_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_305_1 = {2'd0, _zz_when_ArraySlice_l165_305_2};
  assign _zz_when_ArraySlice_l166_305 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_305_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_305_2);
  assign _zz_when_ArraySlice_l166_305_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_305_3);
  assign _zz_when_ArraySlice_l166_305_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_305_3 = {2'd0, _zz_when_ArraySlice_l166_305_4};
  assign _zz__zz_when_ArraySlice_l112_305 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_305 = (_zz_when_ArraySlice_l113_305_1 - _zz_when_ArraySlice_l113_305_4);
  assign _zz_when_ArraySlice_l113_305_1 = (_zz_when_ArraySlice_l113_305_2 + _zz_when_ArraySlice_l113_305_3);
  assign _zz_when_ArraySlice_l113_305_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_305_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_305_4 = {1'd0, _zz_when_ArraySlice_l112_305};
  assign _zz__zz_when_ArraySlice_l173_305 = (_zz__zz_when_ArraySlice_l173_305_1 + _zz__zz_when_ArraySlice_l173_305_2);
  assign _zz__zz_when_ArraySlice_l173_305_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_305_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_305_3 = {1'd0, _zz_when_ArraySlice_l112_305};
  assign _zz_when_ArraySlice_l118_305_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_305 = _zz_when_ArraySlice_l118_305_1[5:0];
  assign _zz_when_ArraySlice_l173_305_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_305_1 = {1'd0, _zz_when_ArraySlice_l173_305_2};
  assign _zz_when_ArraySlice_l173_305_3 = (_zz_when_ArraySlice_l173_305_4 + _zz_when_ArraySlice_l173_305_9);
  assign _zz_when_ArraySlice_l173_305_4 = (_zz_when_ArraySlice_l173_305 - _zz_when_ArraySlice_l173_305_5);
  assign _zz_when_ArraySlice_l173_305_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_305_7);
  assign _zz_when_ArraySlice_l173_305_5 = {1'd0, _zz_when_ArraySlice_l173_305_6};
  assign _zz_when_ArraySlice_l173_305_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_305_7 = {2'd0, _zz_when_ArraySlice_l173_305_8};
  assign _zz_when_ArraySlice_l173_305_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_306 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_306_1);
  assign _zz_when_ArraySlice_l165_306_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_306_1 = {1'd0, _zz_when_ArraySlice_l165_306_2};
  assign _zz_when_ArraySlice_l166_306 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_306_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_306_2);
  assign _zz_when_ArraySlice_l166_306_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_306_3);
  assign _zz_when_ArraySlice_l166_306_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_306_3 = {1'd0, _zz_when_ArraySlice_l166_306_4};
  assign _zz__zz_when_ArraySlice_l112_306 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_306 = (_zz_when_ArraySlice_l113_306_1 - _zz_when_ArraySlice_l113_306_4);
  assign _zz_when_ArraySlice_l113_306_1 = (_zz_when_ArraySlice_l113_306_2 + _zz_when_ArraySlice_l113_306_3);
  assign _zz_when_ArraySlice_l113_306_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_306_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_306_4 = {1'd0, _zz_when_ArraySlice_l112_306};
  assign _zz__zz_when_ArraySlice_l173_306 = (_zz__zz_when_ArraySlice_l173_306_1 + _zz__zz_when_ArraySlice_l173_306_2);
  assign _zz__zz_when_ArraySlice_l173_306_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_306_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_306_3 = {1'd0, _zz_when_ArraySlice_l112_306};
  assign _zz_when_ArraySlice_l118_306_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_306 = _zz_when_ArraySlice_l118_306_1[5:0];
  assign _zz_when_ArraySlice_l173_306_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_306_1 = {1'd0, _zz_when_ArraySlice_l173_306_2};
  assign _zz_when_ArraySlice_l173_306_3 = (_zz_when_ArraySlice_l173_306_4 + _zz_when_ArraySlice_l173_306_9);
  assign _zz_when_ArraySlice_l173_306_4 = (_zz_when_ArraySlice_l173_306 - _zz_when_ArraySlice_l173_306_5);
  assign _zz_when_ArraySlice_l173_306_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_306_7);
  assign _zz_when_ArraySlice_l173_306_5 = {1'd0, _zz_when_ArraySlice_l173_306_6};
  assign _zz_when_ArraySlice_l173_306_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_306_7 = {1'd0, _zz_when_ArraySlice_l173_306_8};
  assign _zz_when_ArraySlice_l173_306_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_307 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_307_1);
  assign _zz_when_ArraySlice_l165_307_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_307_1 = {1'd0, _zz_when_ArraySlice_l165_307_2};
  assign _zz_when_ArraySlice_l166_307 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_307_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_307_2);
  assign _zz_when_ArraySlice_l166_307_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_307_3);
  assign _zz_when_ArraySlice_l166_307_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_307_3 = {1'd0, _zz_when_ArraySlice_l166_307_4};
  assign _zz__zz_when_ArraySlice_l112_307 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_307 = (_zz_when_ArraySlice_l113_307_1 - _zz_when_ArraySlice_l113_307_4);
  assign _zz_when_ArraySlice_l113_307_1 = (_zz_when_ArraySlice_l113_307_2 + _zz_when_ArraySlice_l113_307_3);
  assign _zz_when_ArraySlice_l113_307_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_307_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_307_4 = {1'd0, _zz_when_ArraySlice_l112_307};
  assign _zz__zz_when_ArraySlice_l173_307 = (_zz__zz_when_ArraySlice_l173_307_1 + _zz__zz_when_ArraySlice_l173_307_2);
  assign _zz__zz_when_ArraySlice_l173_307_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_307_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_307_3 = {1'd0, _zz_when_ArraySlice_l112_307};
  assign _zz_when_ArraySlice_l118_307_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_307 = _zz_when_ArraySlice_l118_307_1[5:0];
  assign _zz_when_ArraySlice_l173_307_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_307_1 = {1'd0, _zz_when_ArraySlice_l173_307_2};
  assign _zz_when_ArraySlice_l173_307_3 = (_zz_when_ArraySlice_l173_307_4 + _zz_when_ArraySlice_l173_307_9);
  assign _zz_when_ArraySlice_l173_307_4 = (_zz_when_ArraySlice_l173_307 - _zz_when_ArraySlice_l173_307_5);
  assign _zz_when_ArraySlice_l173_307_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_307_7);
  assign _zz_when_ArraySlice_l173_307_5 = {1'd0, _zz_when_ArraySlice_l173_307_6};
  assign _zz_when_ArraySlice_l173_307_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_307_7 = {1'd0, _zz_when_ArraySlice_l173_307_8};
  assign _zz_when_ArraySlice_l173_307_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_308 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_308_1);
  assign _zz_when_ArraySlice_l165_308_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_308 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_308_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_308_2);
  assign _zz_when_ArraySlice_l166_308_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_308_3);
  assign _zz_when_ArraySlice_l166_308_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_308 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_308 = (_zz_when_ArraySlice_l113_308_1 - _zz_when_ArraySlice_l113_308_4);
  assign _zz_when_ArraySlice_l113_308_1 = (_zz_when_ArraySlice_l113_308_2 + _zz_when_ArraySlice_l113_308_3);
  assign _zz_when_ArraySlice_l113_308_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_308_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_308_4 = {1'd0, _zz_when_ArraySlice_l112_308};
  assign _zz__zz_when_ArraySlice_l173_308 = (_zz__zz_when_ArraySlice_l173_308_1 + _zz__zz_when_ArraySlice_l173_308_2);
  assign _zz__zz_when_ArraySlice_l173_308_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_308_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_308_3 = {1'd0, _zz_when_ArraySlice_l112_308};
  assign _zz_when_ArraySlice_l118_308_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_308 = _zz_when_ArraySlice_l118_308_1[5:0];
  assign _zz_when_ArraySlice_l173_308_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_308_1 = {1'd0, _zz_when_ArraySlice_l173_308_2};
  assign _zz_when_ArraySlice_l173_308_3 = (_zz_when_ArraySlice_l173_308_4 + _zz_when_ArraySlice_l173_308_8);
  assign _zz_when_ArraySlice_l173_308_4 = (_zz_when_ArraySlice_l173_308 - _zz_when_ArraySlice_l173_308_5);
  assign _zz_when_ArraySlice_l173_308_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_308_7);
  assign _zz_when_ArraySlice_l173_308_5 = {1'd0, _zz_when_ArraySlice_l173_308_6};
  assign _zz_when_ArraySlice_l173_308_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_308_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_309 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_309_1);
  assign _zz_when_ArraySlice_l165_309_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_309_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_309 = {1'd0, _zz_when_ArraySlice_l166_309_1};
  assign _zz_when_ArraySlice_l166_309_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_309_3);
  assign _zz_when_ArraySlice_l166_309_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_309_4);
  assign _zz_when_ArraySlice_l166_309_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_309 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_309 = (_zz_when_ArraySlice_l113_309_1 - _zz_when_ArraySlice_l113_309_4);
  assign _zz_when_ArraySlice_l113_309_1 = (_zz_when_ArraySlice_l113_309_2 + _zz_when_ArraySlice_l113_309_3);
  assign _zz_when_ArraySlice_l113_309_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_309_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_309_4 = {1'd0, _zz_when_ArraySlice_l112_309};
  assign _zz__zz_when_ArraySlice_l173_309 = (_zz__zz_when_ArraySlice_l173_309_1 + _zz__zz_when_ArraySlice_l173_309_2);
  assign _zz__zz_when_ArraySlice_l173_309_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_309_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_309_3 = {1'd0, _zz_when_ArraySlice_l112_309};
  assign _zz_when_ArraySlice_l118_309_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_309 = _zz_when_ArraySlice_l118_309_1[5:0];
  assign _zz_when_ArraySlice_l173_309_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_309_1 = {2'd0, _zz_when_ArraySlice_l173_309_2};
  assign _zz_when_ArraySlice_l173_309_3 = (_zz_when_ArraySlice_l173_309_4 + _zz_when_ArraySlice_l173_309_8);
  assign _zz_when_ArraySlice_l173_309_4 = (_zz_when_ArraySlice_l173_309 - _zz_when_ArraySlice_l173_309_5);
  assign _zz_when_ArraySlice_l173_309_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_309_7);
  assign _zz_when_ArraySlice_l173_309_5 = {1'd0, _zz_when_ArraySlice_l173_309_6};
  assign _zz_when_ArraySlice_l173_309_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_309_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_310 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_310_1);
  assign _zz_when_ArraySlice_l165_310_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_310_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_310 = {1'd0, _zz_when_ArraySlice_l166_310_1};
  assign _zz_when_ArraySlice_l166_310_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_310_3);
  assign _zz_when_ArraySlice_l166_310_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_310_4);
  assign _zz_when_ArraySlice_l166_310_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_310 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_310 = (_zz_when_ArraySlice_l113_310_1 - _zz_when_ArraySlice_l113_310_4);
  assign _zz_when_ArraySlice_l113_310_1 = (_zz_when_ArraySlice_l113_310_2 + _zz_when_ArraySlice_l113_310_3);
  assign _zz_when_ArraySlice_l113_310_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_310_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_310_4 = {1'd0, _zz_when_ArraySlice_l112_310};
  assign _zz__zz_when_ArraySlice_l173_310 = (_zz__zz_when_ArraySlice_l173_310_1 + _zz__zz_when_ArraySlice_l173_310_2);
  assign _zz__zz_when_ArraySlice_l173_310_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_310_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_310_3 = {1'd0, _zz_when_ArraySlice_l112_310};
  assign _zz_when_ArraySlice_l118_310_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_310 = _zz_when_ArraySlice_l118_310_1[5:0];
  assign _zz_when_ArraySlice_l173_310_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_310_1 = {2'd0, _zz_when_ArraySlice_l173_310_2};
  assign _zz_when_ArraySlice_l173_310_3 = (_zz_when_ArraySlice_l173_310_4 + _zz_when_ArraySlice_l173_310_8);
  assign _zz_when_ArraySlice_l173_310_4 = (_zz_when_ArraySlice_l173_310 - _zz_when_ArraySlice_l173_310_5);
  assign _zz_when_ArraySlice_l173_310_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_310_7);
  assign _zz_when_ArraySlice_l173_310_5 = {1'd0, _zz_when_ArraySlice_l173_310_6};
  assign _zz_when_ArraySlice_l173_310_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_310_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_311 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_311_1);
  assign _zz_when_ArraySlice_l165_311_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_311_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_311 = {2'd0, _zz_when_ArraySlice_l166_311_1};
  assign _zz_when_ArraySlice_l166_311_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_311_3);
  assign _zz_when_ArraySlice_l166_311_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_311_4);
  assign _zz_when_ArraySlice_l166_311_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_311 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_311 = (_zz_when_ArraySlice_l113_311_1 - _zz_when_ArraySlice_l113_311_4);
  assign _zz_when_ArraySlice_l113_311_1 = (_zz_when_ArraySlice_l113_311_2 + _zz_when_ArraySlice_l113_311_3);
  assign _zz_when_ArraySlice_l113_311_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_311_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_311_4 = {1'd0, _zz_when_ArraySlice_l112_311};
  assign _zz__zz_when_ArraySlice_l173_311 = (_zz__zz_when_ArraySlice_l173_311_1 + _zz__zz_when_ArraySlice_l173_311_2);
  assign _zz__zz_when_ArraySlice_l173_311_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_311_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_311_3 = {1'd0, _zz_when_ArraySlice_l112_311};
  assign _zz_when_ArraySlice_l118_311_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_311 = _zz_when_ArraySlice_l118_311_1[5:0];
  assign _zz_when_ArraySlice_l173_311_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_311_1 = {3'd0, _zz_when_ArraySlice_l173_311_2};
  assign _zz_when_ArraySlice_l173_311_3 = (_zz_when_ArraySlice_l173_311_4 + _zz_when_ArraySlice_l173_311_8);
  assign _zz_when_ArraySlice_l173_311_4 = (_zz_when_ArraySlice_l173_311 - _zz_when_ArraySlice_l173_311_5);
  assign _zz_when_ArraySlice_l173_311_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_311_7);
  assign _zz_when_ArraySlice_l173_311_5 = {1'd0, _zz_when_ArraySlice_l173_311_6};
  assign _zz_when_ArraySlice_l173_311_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_311_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l268_4_1 = (_zz_when_ArraySlice_l268_4_2 + _zz_when_ArraySlice_l268_4_7);
  assign _zz_when_ArraySlice_l268_4_2 = (_zz_when_ArraySlice_l268_4_3 + _zz_when_ArraySlice_l268_4_5);
  assign _zz_when_ArraySlice_l268_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l268_4_4);
  assign _zz_when_ArraySlice_l268_4_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l268_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l268_4_5 = {5'd0, _zz_when_ArraySlice_l268_4_6};
  assign _zz_when_ArraySlice_l268_4_7 = (bReg * 3'b100);
  assign _zz_selectReadFifo_4_47 = 1'b1;
  assign _zz_selectReadFifo_4_46 = {5'd0, _zz_selectReadFifo_4_47};
  assign _zz_when_ArraySlice_l272_4 = (_zz_when_ArraySlice_l272_4_1 % aReg);
  assign _zz_when_ArraySlice_l272_4_1 = (handshakeTimes_4_value + _zz_when_ArraySlice_l272_4_2);
  assign _zz_when_ArraySlice_l272_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l272_4_2 = {12'd0, _zz_when_ArraySlice_l272_4_3};
  assign _zz_when_ArraySlice_l276_4_1 = (selectReadFifo_4 + _zz_when_ArraySlice_l276_4_2);
  assign _zz_when_ArraySlice_l276_4_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l277_4_2 = (_zz_when_ArraySlice_l277_4_3 - _zz_when_ArraySlice_l277_4_4);
  assign _zz_when_ArraySlice_l277_4_1 = {7'd0, _zz_when_ArraySlice_l277_4_2};
  assign _zz_when_ArraySlice_l277_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l277_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l277_4_4 = {5'd0, _zz_when_ArraySlice_l277_4_5};
  assign _zz__zz_when_ArraySlice_l94_37 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_37 = (_zz_when_ArraySlice_l95_37_1 - _zz_when_ArraySlice_l95_37_4);
  assign _zz_when_ArraySlice_l95_37_1 = (_zz_when_ArraySlice_l95_37_2 + _zz_when_ArraySlice_l95_37_3);
  assign _zz_when_ArraySlice_l95_37_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_37_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_37_4 = {1'd0, _zz_when_ArraySlice_l94_37};
  assign _zz__zz_when_ArraySlice_l279_4 = (_zz__zz_when_ArraySlice_l279_4_1 + _zz__zz_when_ArraySlice_l279_4_2);
  assign _zz__zz_when_ArraySlice_l279_4_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l279_4_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l279_4_3 = {1'd0, _zz_when_ArraySlice_l94_37};
  assign _zz_when_ArraySlice_l99_37_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_37 = _zz_when_ArraySlice_l99_37_1[5:0];
  assign _zz_when_ArraySlice_l279_4_1 = (outSliceNumb_4_value + _zz_when_ArraySlice_l279_4_2);
  assign _zz_when_ArraySlice_l279_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l279_4_2 = {6'd0, _zz_when_ArraySlice_l279_4_3};
  assign _zz_when_ArraySlice_l279_4_4 = (_zz_when_ArraySlice_l279_4 / aReg);
  assign _zz_selectReadFifo_4_48 = (selectReadFifo_4 - _zz_selectReadFifo_4_49);
  assign _zz_selectReadFifo_4_49 = {3'd0, bReg};
  assign _zz_selectReadFifo_4_51 = 1'b1;
  assign _zz_selectReadFifo_4_50 = {5'd0, _zz_selectReadFifo_4_51};
  assign _zz_selectReadFifo_4_52 = (selectReadFifo_4 + _zz_selectReadFifo_4_53);
  assign _zz_selectReadFifo_4_53 = (3'b111 * bReg);
  assign _zz_selectReadFifo_4_55 = 1'b1;
  assign _zz_selectReadFifo_4_54 = {5'd0, _zz_selectReadFifo_4_55};
  assign _zz_when_ArraySlice_l165_312 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_312_1);
  assign _zz_when_ArraySlice_l165_312_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_312_1 = {3'd0, _zz_when_ArraySlice_l165_312_2};
  assign _zz_when_ArraySlice_l166_312 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_312_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_312_3);
  assign _zz_when_ArraySlice_l166_312_1 = {1'd0, _zz_when_ArraySlice_l166_312_2};
  assign _zz_when_ArraySlice_l166_312_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_312_4);
  assign _zz_when_ArraySlice_l166_312_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_312_4 = {3'd0, _zz_when_ArraySlice_l166_312_5};
  assign _zz__zz_when_ArraySlice_l112_312 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_312 = (_zz_when_ArraySlice_l113_312_1 - _zz_when_ArraySlice_l113_312_4);
  assign _zz_when_ArraySlice_l113_312_1 = (_zz_when_ArraySlice_l113_312_2 + _zz_when_ArraySlice_l113_312_3);
  assign _zz_when_ArraySlice_l113_312_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_312_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_312_4 = {1'd0, _zz_when_ArraySlice_l112_312};
  assign _zz__zz_when_ArraySlice_l173_312 = (_zz__zz_when_ArraySlice_l173_312_1 + _zz__zz_when_ArraySlice_l173_312_2);
  assign _zz__zz_when_ArraySlice_l173_312_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_312_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_312_3 = {1'd0, _zz_when_ArraySlice_l112_312};
  assign _zz_when_ArraySlice_l118_312_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_312 = _zz_when_ArraySlice_l118_312_1[5:0];
  assign _zz_when_ArraySlice_l173_312_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_312_2 = (_zz_when_ArraySlice_l173_312_3 + _zz_when_ArraySlice_l173_312_8);
  assign _zz_when_ArraySlice_l173_312_3 = (_zz_when_ArraySlice_l173_312 - _zz_when_ArraySlice_l173_312_4);
  assign _zz_when_ArraySlice_l173_312_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_312_6);
  assign _zz_when_ArraySlice_l173_312_4 = {1'd0, _zz_when_ArraySlice_l173_312_5};
  assign _zz_when_ArraySlice_l173_312_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_312_6 = {3'd0, _zz_when_ArraySlice_l173_312_7};
  assign _zz_when_ArraySlice_l173_312_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_313 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_313_1);
  assign _zz_when_ArraySlice_l165_313_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_313_1 = {2'd0, _zz_when_ArraySlice_l165_313_2};
  assign _zz_when_ArraySlice_l166_313 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_313_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_313_2);
  assign _zz_when_ArraySlice_l166_313_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_313_3);
  assign _zz_when_ArraySlice_l166_313_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_313_3 = {2'd0, _zz_when_ArraySlice_l166_313_4};
  assign _zz__zz_when_ArraySlice_l112_313 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_313 = (_zz_when_ArraySlice_l113_313_1 - _zz_when_ArraySlice_l113_313_4);
  assign _zz_when_ArraySlice_l113_313_1 = (_zz_when_ArraySlice_l113_313_2 + _zz_when_ArraySlice_l113_313_3);
  assign _zz_when_ArraySlice_l113_313_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_313_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_313_4 = {1'd0, _zz_when_ArraySlice_l112_313};
  assign _zz__zz_when_ArraySlice_l173_313 = (_zz__zz_when_ArraySlice_l173_313_1 + _zz__zz_when_ArraySlice_l173_313_2);
  assign _zz__zz_when_ArraySlice_l173_313_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_313_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_313_3 = {1'd0, _zz_when_ArraySlice_l112_313};
  assign _zz_when_ArraySlice_l118_313_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_313 = _zz_when_ArraySlice_l118_313_1[5:0];
  assign _zz_when_ArraySlice_l173_313_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_313_1 = {1'd0, _zz_when_ArraySlice_l173_313_2};
  assign _zz_when_ArraySlice_l173_313_3 = (_zz_when_ArraySlice_l173_313_4 + _zz_when_ArraySlice_l173_313_9);
  assign _zz_when_ArraySlice_l173_313_4 = (_zz_when_ArraySlice_l173_313 - _zz_when_ArraySlice_l173_313_5);
  assign _zz_when_ArraySlice_l173_313_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_313_7);
  assign _zz_when_ArraySlice_l173_313_5 = {1'd0, _zz_when_ArraySlice_l173_313_6};
  assign _zz_when_ArraySlice_l173_313_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_313_7 = {2'd0, _zz_when_ArraySlice_l173_313_8};
  assign _zz_when_ArraySlice_l173_313_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_314 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_314_1);
  assign _zz_when_ArraySlice_l165_314_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_314_1 = {1'd0, _zz_when_ArraySlice_l165_314_2};
  assign _zz_when_ArraySlice_l166_314 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_314_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_314_2);
  assign _zz_when_ArraySlice_l166_314_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_314_3);
  assign _zz_when_ArraySlice_l166_314_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_314_3 = {1'd0, _zz_when_ArraySlice_l166_314_4};
  assign _zz__zz_when_ArraySlice_l112_314 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_314 = (_zz_when_ArraySlice_l113_314_1 - _zz_when_ArraySlice_l113_314_4);
  assign _zz_when_ArraySlice_l113_314_1 = (_zz_when_ArraySlice_l113_314_2 + _zz_when_ArraySlice_l113_314_3);
  assign _zz_when_ArraySlice_l113_314_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_314_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_314_4 = {1'd0, _zz_when_ArraySlice_l112_314};
  assign _zz__zz_when_ArraySlice_l173_314 = (_zz__zz_when_ArraySlice_l173_314_1 + _zz__zz_when_ArraySlice_l173_314_2);
  assign _zz__zz_when_ArraySlice_l173_314_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_314_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_314_3 = {1'd0, _zz_when_ArraySlice_l112_314};
  assign _zz_when_ArraySlice_l118_314_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_314 = _zz_when_ArraySlice_l118_314_1[5:0];
  assign _zz_when_ArraySlice_l173_314_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_314_1 = {1'd0, _zz_when_ArraySlice_l173_314_2};
  assign _zz_when_ArraySlice_l173_314_3 = (_zz_when_ArraySlice_l173_314_4 + _zz_when_ArraySlice_l173_314_9);
  assign _zz_when_ArraySlice_l173_314_4 = (_zz_when_ArraySlice_l173_314 - _zz_when_ArraySlice_l173_314_5);
  assign _zz_when_ArraySlice_l173_314_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_314_7);
  assign _zz_when_ArraySlice_l173_314_5 = {1'd0, _zz_when_ArraySlice_l173_314_6};
  assign _zz_when_ArraySlice_l173_314_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_314_7 = {1'd0, _zz_when_ArraySlice_l173_314_8};
  assign _zz_when_ArraySlice_l173_314_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_315 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_315_1);
  assign _zz_when_ArraySlice_l165_315_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_315_1 = {1'd0, _zz_when_ArraySlice_l165_315_2};
  assign _zz_when_ArraySlice_l166_315 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_315_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_315_2);
  assign _zz_when_ArraySlice_l166_315_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_315_3);
  assign _zz_when_ArraySlice_l166_315_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_315_3 = {1'd0, _zz_when_ArraySlice_l166_315_4};
  assign _zz__zz_when_ArraySlice_l112_315 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_315 = (_zz_when_ArraySlice_l113_315_1 - _zz_when_ArraySlice_l113_315_4);
  assign _zz_when_ArraySlice_l113_315_1 = (_zz_when_ArraySlice_l113_315_2 + _zz_when_ArraySlice_l113_315_3);
  assign _zz_when_ArraySlice_l113_315_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_315_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_315_4 = {1'd0, _zz_when_ArraySlice_l112_315};
  assign _zz__zz_when_ArraySlice_l173_315 = (_zz__zz_when_ArraySlice_l173_315_1 + _zz__zz_when_ArraySlice_l173_315_2);
  assign _zz__zz_when_ArraySlice_l173_315_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_315_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_315_3 = {1'd0, _zz_when_ArraySlice_l112_315};
  assign _zz_when_ArraySlice_l118_315_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_315 = _zz_when_ArraySlice_l118_315_1[5:0];
  assign _zz_when_ArraySlice_l173_315_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_315_1 = {1'd0, _zz_when_ArraySlice_l173_315_2};
  assign _zz_when_ArraySlice_l173_315_3 = (_zz_when_ArraySlice_l173_315_4 + _zz_when_ArraySlice_l173_315_9);
  assign _zz_when_ArraySlice_l173_315_4 = (_zz_when_ArraySlice_l173_315 - _zz_when_ArraySlice_l173_315_5);
  assign _zz_when_ArraySlice_l173_315_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_315_7);
  assign _zz_when_ArraySlice_l173_315_5 = {1'd0, _zz_when_ArraySlice_l173_315_6};
  assign _zz_when_ArraySlice_l173_315_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_315_7 = {1'd0, _zz_when_ArraySlice_l173_315_8};
  assign _zz_when_ArraySlice_l173_315_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_316 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_316_1);
  assign _zz_when_ArraySlice_l165_316_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_316 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_316_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_316_2);
  assign _zz_when_ArraySlice_l166_316_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_316_3);
  assign _zz_when_ArraySlice_l166_316_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_316 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_316 = (_zz_when_ArraySlice_l113_316_1 - _zz_when_ArraySlice_l113_316_4);
  assign _zz_when_ArraySlice_l113_316_1 = (_zz_when_ArraySlice_l113_316_2 + _zz_when_ArraySlice_l113_316_3);
  assign _zz_when_ArraySlice_l113_316_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_316_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_316_4 = {1'd0, _zz_when_ArraySlice_l112_316};
  assign _zz__zz_when_ArraySlice_l173_316 = (_zz__zz_when_ArraySlice_l173_316_1 + _zz__zz_when_ArraySlice_l173_316_2);
  assign _zz__zz_when_ArraySlice_l173_316_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_316_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_316_3 = {1'd0, _zz_when_ArraySlice_l112_316};
  assign _zz_when_ArraySlice_l118_316_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_316 = _zz_when_ArraySlice_l118_316_1[5:0];
  assign _zz_when_ArraySlice_l173_316_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_316_1 = {1'd0, _zz_when_ArraySlice_l173_316_2};
  assign _zz_when_ArraySlice_l173_316_3 = (_zz_when_ArraySlice_l173_316_4 + _zz_when_ArraySlice_l173_316_8);
  assign _zz_when_ArraySlice_l173_316_4 = (_zz_when_ArraySlice_l173_316 - _zz_when_ArraySlice_l173_316_5);
  assign _zz_when_ArraySlice_l173_316_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_316_7);
  assign _zz_when_ArraySlice_l173_316_5 = {1'd0, _zz_when_ArraySlice_l173_316_6};
  assign _zz_when_ArraySlice_l173_316_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_316_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_317 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_317_1);
  assign _zz_when_ArraySlice_l165_317_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_317_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_317 = {1'd0, _zz_when_ArraySlice_l166_317_1};
  assign _zz_when_ArraySlice_l166_317_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_317_3);
  assign _zz_when_ArraySlice_l166_317_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_317_4);
  assign _zz_when_ArraySlice_l166_317_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_317 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_317 = (_zz_when_ArraySlice_l113_317_1 - _zz_when_ArraySlice_l113_317_4);
  assign _zz_when_ArraySlice_l113_317_1 = (_zz_when_ArraySlice_l113_317_2 + _zz_when_ArraySlice_l113_317_3);
  assign _zz_when_ArraySlice_l113_317_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_317_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_317_4 = {1'd0, _zz_when_ArraySlice_l112_317};
  assign _zz__zz_when_ArraySlice_l173_317 = (_zz__zz_when_ArraySlice_l173_317_1 + _zz__zz_when_ArraySlice_l173_317_2);
  assign _zz__zz_when_ArraySlice_l173_317_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_317_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_317_3 = {1'd0, _zz_when_ArraySlice_l112_317};
  assign _zz_when_ArraySlice_l118_317_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_317 = _zz_when_ArraySlice_l118_317_1[5:0];
  assign _zz_when_ArraySlice_l173_317_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_317_1 = {2'd0, _zz_when_ArraySlice_l173_317_2};
  assign _zz_when_ArraySlice_l173_317_3 = (_zz_when_ArraySlice_l173_317_4 + _zz_when_ArraySlice_l173_317_8);
  assign _zz_when_ArraySlice_l173_317_4 = (_zz_when_ArraySlice_l173_317 - _zz_when_ArraySlice_l173_317_5);
  assign _zz_when_ArraySlice_l173_317_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_317_7);
  assign _zz_when_ArraySlice_l173_317_5 = {1'd0, _zz_when_ArraySlice_l173_317_6};
  assign _zz_when_ArraySlice_l173_317_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_317_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_318 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_318_1);
  assign _zz_when_ArraySlice_l165_318_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_318_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_318 = {1'd0, _zz_when_ArraySlice_l166_318_1};
  assign _zz_when_ArraySlice_l166_318_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_318_3);
  assign _zz_when_ArraySlice_l166_318_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_318_4);
  assign _zz_when_ArraySlice_l166_318_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_318 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_318 = (_zz_when_ArraySlice_l113_318_1 - _zz_when_ArraySlice_l113_318_4);
  assign _zz_when_ArraySlice_l113_318_1 = (_zz_when_ArraySlice_l113_318_2 + _zz_when_ArraySlice_l113_318_3);
  assign _zz_when_ArraySlice_l113_318_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_318_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_318_4 = {1'd0, _zz_when_ArraySlice_l112_318};
  assign _zz__zz_when_ArraySlice_l173_318 = (_zz__zz_when_ArraySlice_l173_318_1 + _zz__zz_when_ArraySlice_l173_318_2);
  assign _zz__zz_when_ArraySlice_l173_318_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_318_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_318_3 = {1'd0, _zz_when_ArraySlice_l112_318};
  assign _zz_when_ArraySlice_l118_318_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_318 = _zz_when_ArraySlice_l118_318_1[5:0];
  assign _zz_when_ArraySlice_l173_318_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_318_1 = {2'd0, _zz_when_ArraySlice_l173_318_2};
  assign _zz_when_ArraySlice_l173_318_3 = (_zz_when_ArraySlice_l173_318_4 + _zz_when_ArraySlice_l173_318_8);
  assign _zz_when_ArraySlice_l173_318_4 = (_zz_when_ArraySlice_l173_318 - _zz_when_ArraySlice_l173_318_5);
  assign _zz_when_ArraySlice_l173_318_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_318_7);
  assign _zz_when_ArraySlice_l173_318_5 = {1'd0, _zz_when_ArraySlice_l173_318_6};
  assign _zz_when_ArraySlice_l173_318_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_318_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_319 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_319_1);
  assign _zz_when_ArraySlice_l165_319_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_319_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_319 = {2'd0, _zz_when_ArraySlice_l166_319_1};
  assign _zz_when_ArraySlice_l166_319_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_319_3);
  assign _zz_when_ArraySlice_l166_319_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_319_4);
  assign _zz_when_ArraySlice_l166_319_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_319 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_319 = (_zz_when_ArraySlice_l113_319_1 - _zz_when_ArraySlice_l113_319_4);
  assign _zz_when_ArraySlice_l113_319_1 = (_zz_when_ArraySlice_l113_319_2 + _zz_when_ArraySlice_l113_319_3);
  assign _zz_when_ArraySlice_l113_319_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_319_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_319_4 = {1'd0, _zz_when_ArraySlice_l112_319};
  assign _zz__zz_when_ArraySlice_l173_319 = (_zz__zz_when_ArraySlice_l173_319_1 + _zz__zz_when_ArraySlice_l173_319_2);
  assign _zz__zz_when_ArraySlice_l173_319_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_319_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_319_3 = {1'd0, _zz_when_ArraySlice_l112_319};
  assign _zz_when_ArraySlice_l118_319_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_319 = _zz_when_ArraySlice_l118_319_1[5:0];
  assign _zz_when_ArraySlice_l173_319_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_319_1 = {3'd0, _zz_when_ArraySlice_l173_319_2};
  assign _zz_when_ArraySlice_l173_319_3 = (_zz_when_ArraySlice_l173_319_4 + _zz_when_ArraySlice_l173_319_8);
  assign _zz_when_ArraySlice_l173_319_4 = (_zz_when_ArraySlice_l173_319 - _zz_when_ArraySlice_l173_319_5);
  assign _zz_when_ArraySlice_l173_319_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_319_7);
  assign _zz_when_ArraySlice_l173_319_5 = {1'd0, _zz_when_ArraySlice_l173_319_6};
  assign _zz_when_ArraySlice_l173_319_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_319_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l288_4_1 = (_zz_when_ArraySlice_l288_4_2 + _zz_when_ArraySlice_l288_4_7);
  assign _zz_when_ArraySlice_l288_4_2 = (_zz_when_ArraySlice_l288_4_3 + _zz_when_ArraySlice_l288_4_5);
  assign _zz_when_ArraySlice_l288_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l288_4_4);
  assign _zz_when_ArraySlice_l288_4_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l288_4_5 = {5'd0, _zz_when_ArraySlice_l288_4_6};
  assign _zz_when_ArraySlice_l288_4_7 = (bReg * 3'b100);
  assign _zz_selectReadFifo_4_57 = 1'b1;
  assign _zz_selectReadFifo_4_56 = {5'd0, _zz_selectReadFifo_4_57};
  assign _zz_when_ArraySlice_l292_4 = (_zz_when_ArraySlice_l292_4_1 % aReg);
  assign _zz_when_ArraySlice_l292_4_1 = (handshakeTimes_4_value + _zz_when_ArraySlice_l292_4_2);
  assign _zz_when_ArraySlice_l292_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l292_4_2 = {12'd0, _zz_when_ArraySlice_l292_4_3};
  assign _zz_when_ArraySlice_l303_4_2 = (_zz_when_ArraySlice_l303_4_3 - _zz_when_ArraySlice_l303_4_4);
  assign _zz_when_ArraySlice_l303_4_1 = {7'd0, _zz_when_ArraySlice_l303_4_2};
  assign _zz_when_ArraySlice_l303_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l303_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l303_4_4 = {5'd0, _zz_when_ArraySlice_l303_4_5};
  assign _zz__zz_when_ArraySlice_l94_38 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_38 = (_zz_when_ArraySlice_l95_38_1 - _zz_when_ArraySlice_l95_38_4);
  assign _zz_when_ArraySlice_l95_38_1 = (_zz_when_ArraySlice_l95_38_2 + _zz_when_ArraySlice_l95_38_3);
  assign _zz_when_ArraySlice_l95_38_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_38_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_38_4 = {1'd0, _zz_when_ArraySlice_l94_38};
  assign _zz__zz_when_ArraySlice_l304_4 = (_zz__zz_when_ArraySlice_l304_4_1 + _zz__zz_when_ArraySlice_l304_4_2);
  assign _zz__zz_when_ArraySlice_l304_4_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l304_4_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l304_4_3 = {1'd0, _zz_when_ArraySlice_l94_38};
  assign _zz_when_ArraySlice_l99_38_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_38 = _zz_when_ArraySlice_l99_38_1[5:0];
  assign _zz_when_ArraySlice_l304_4_1 = (outSliceNumb_4_value + _zz_when_ArraySlice_l304_4_2);
  assign _zz_when_ArraySlice_l304_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l304_4_2 = {6'd0, _zz_when_ArraySlice_l304_4_3};
  assign _zz_when_ArraySlice_l304_4_4 = (_zz_when_ArraySlice_l304_4 / aReg);
  assign _zz_selectReadFifo_4_58 = (selectReadFifo_4 - _zz_selectReadFifo_4_59);
  assign _zz_selectReadFifo_4_59 = {3'd0, bReg};
  assign _zz_selectReadFifo_4_61 = 1'b1;
  assign _zz_selectReadFifo_4_60 = {5'd0, _zz_selectReadFifo_4_61};
  assign _zz_when_ArraySlice_l165_320 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_320_1);
  assign _zz_when_ArraySlice_l165_320_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_320_1 = {3'd0, _zz_when_ArraySlice_l165_320_2};
  assign _zz_when_ArraySlice_l166_320 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_320_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_320_3);
  assign _zz_when_ArraySlice_l166_320_1 = {1'd0, _zz_when_ArraySlice_l166_320_2};
  assign _zz_when_ArraySlice_l166_320_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_320_4);
  assign _zz_when_ArraySlice_l166_320_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_320_4 = {3'd0, _zz_when_ArraySlice_l166_320_5};
  assign _zz__zz_when_ArraySlice_l112_320 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_320 = (_zz_when_ArraySlice_l113_320_1 - _zz_when_ArraySlice_l113_320_4);
  assign _zz_when_ArraySlice_l113_320_1 = (_zz_when_ArraySlice_l113_320_2 + _zz_when_ArraySlice_l113_320_3);
  assign _zz_when_ArraySlice_l113_320_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_320_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_320_4 = {1'd0, _zz_when_ArraySlice_l112_320};
  assign _zz__zz_when_ArraySlice_l173_320 = (_zz__zz_when_ArraySlice_l173_320_1 + _zz__zz_when_ArraySlice_l173_320_2);
  assign _zz__zz_when_ArraySlice_l173_320_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_320_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_320_3 = {1'd0, _zz_when_ArraySlice_l112_320};
  assign _zz_when_ArraySlice_l118_320_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_320 = _zz_when_ArraySlice_l118_320_1[5:0];
  assign _zz_when_ArraySlice_l173_320_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_320_2 = (_zz_when_ArraySlice_l173_320_3 + _zz_when_ArraySlice_l173_320_8);
  assign _zz_when_ArraySlice_l173_320_3 = (_zz_when_ArraySlice_l173_320 - _zz_when_ArraySlice_l173_320_4);
  assign _zz_when_ArraySlice_l173_320_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_320_6);
  assign _zz_when_ArraySlice_l173_320_4 = {1'd0, _zz_when_ArraySlice_l173_320_5};
  assign _zz_when_ArraySlice_l173_320_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_320_6 = {3'd0, _zz_when_ArraySlice_l173_320_7};
  assign _zz_when_ArraySlice_l173_320_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_321 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_321_1);
  assign _zz_when_ArraySlice_l165_321_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_321_1 = {2'd0, _zz_when_ArraySlice_l165_321_2};
  assign _zz_when_ArraySlice_l166_321 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_321_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_321_2);
  assign _zz_when_ArraySlice_l166_321_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_321_3);
  assign _zz_when_ArraySlice_l166_321_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_321_3 = {2'd0, _zz_when_ArraySlice_l166_321_4};
  assign _zz__zz_when_ArraySlice_l112_321 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_321 = (_zz_when_ArraySlice_l113_321_1 - _zz_when_ArraySlice_l113_321_4);
  assign _zz_when_ArraySlice_l113_321_1 = (_zz_when_ArraySlice_l113_321_2 + _zz_when_ArraySlice_l113_321_3);
  assign _zz_when_ArraySlice_l113_321_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_321_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_321_4 = {1'd0, _zz_when_ArraySlice_l112_321};
  assign _zz__zz_when_ArraySlice_l173_321 = (_zz__zz_when_ArraySlice_l173_321_1 + _zz__zz_when_ArraySlice_l173_321_2);
  assign _zz__zz_when_ArraySlice_l173_321_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_321_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_321_3 = {1'd0, _zz_when_ArraySlice_l112_321};
  assign _zz_when_ArraySlice_l118_321_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_321 = _zz_when_ArraySlice_l118_321_1[5:0];
  assign _zz_when_ArraySlice_l173_321_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_321_1 = {1'd0, _zz_when_ArraySlice_l173_321_2};
  assign _zz_when_ArraySlice_l173_321_3 = (_zz_when_ArraySlice_l173_321_4 + _zz_when_ArraySlice_l173_321_9);
  assign _zz_when_ArraySlice_l173_321_4 = (_zz_when_ArraySlice_l173_321 - _zz_when_ArraySlice_l173_321_5);
  assign _zz_when_ArraySlice_l173_321_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_321_7);
  assign _zz_when_ArraySlice_l173_321_5 = {1'd0, _zz_when_ArraySlice_l173_321_6};
  assign _zz_when_ArraySlice_l173_321_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_321_7 = {2'd0, _zz_when_ArraySlice_l173_321_8};
  assign _zz_when_ArraySlice_l173_321_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_322 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_322_1);
  assign _zz_when_ArraySlice_l165_322_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_322_1 = {1'd0, _zz_when_ArraySlice_l165_322_2};
  assign _zz_when_ArraySlice_l166_322 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_322_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_322_2);
  assign _zz_when_ArraySlice_l166_322_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_322_3);
  assign _zz_when_ArraySlice_l166_322_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_322_3 = {1'd0, _zz_when_ArraySlice_l166_322_4};
  assign _zz__zz_when_ArraySlice_l112_322 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_322 = (_zz_when_ArraySlice_l113_322_1 - _zz_when_ArraySlice_l113_322_4);
  assign _zz_when_ArraySlice_l113_322_1 = (_zz_when_ArraySlice_l113_322_2 + _zz_when_ArraySlice_l113_322_3);
  assign _zz_when_ArraySlice_l113_322_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_322_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_322_4 = {1'd0, _zz_when_ArraySlice_l112_322};
  assign _zz__zz_when_ArraySlice_l173_322 = (_zz__zz_when_ArraySlice_l173_322_1 + _zz__zz_when_ArraySlice_l173_322_2);
  assign _zz__zz_when_ArraySlice_l173_322_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_322_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_322_3 = {1'd0, _zz_when_ArraySlice_l112_322};
  assign _zz_when_ArraySlice_l118_322_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_322 = _zz_when_ArraySlice_l118_322_1[5:0];
  assign _zz_when_ArraySlice_l173_322_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_322_1 = {1'd0, _zz_when_ArraySlice_l173_322_2};
  assign _zz_when_ArraySlice_l173_322_3 = (_zz_when_ArraySlice_l173_322_4 + _zz_when_ArraySlice_l173_322_9);
  assign _zz_when_ArraySlice_l173_322_4 = (_zz_when_ArraySlice_l173_322 - _zz_when_ArraySlice_l173_322_5);
  assign _zz_when_ArraySlice_l173_322_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_322_7);
  assign _zz_when_ArraySlice_l173_322_5 = {1'd0, _zz_when_ArraySlice_l173_322_6};
  assign _zz_when_ArraySlice_l173_322_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_322_7 = {1'd0, _zz_when_ArraySlice_l173_322_8};
  assign _zz_when_ArraySlice_l173_322_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_323 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_323_1);
  assign _zz_when_ArraySlice_l165_323_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_323_1 = {1'd0, _zz_when_ArraySlice_l165_323_2};
  assign _zz_when_ArraySlice_l166_323 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_323_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_323_2);
  assign _zz_when_ArraySlice_l166_323_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_323_3);
  assign _zz_when_ArraySlice_l166_323_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_323_3 = {1'd0, _zz_when_ArraySlice_l166_323_4};
  assign _zz__zz_when_ArraySlice_l112_323 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_323 = (_zz_when_ArraySlice_l113_323_1 - _zz_when_ArraySlice_l113_323_4);
  assign _zz_when_ArraySlice_l113_323_1 = (_zz_when_ArraySlice_l113_323_2 + _zz_when_ArraySlice_l113_323_3);
  assign _zz_when_ArraySlice_l113_323_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_323_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_323_4 = {1'd0, _zz_when_ArraySlice_l112_323};
  assign _zz__zz_when_ArraySlice_l173_323 = (_zz__zz_when_ArraySlice_l173_323_1 + _zz__zz_when_ArraySlice_l173_323_2);
  assign _zz__zz_when_ArraySlice_l173_323_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_323_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_323_3 = {1'd0, _zz_when_ArraySlice_l112_323};
  assign _zz_when_ArraySlice_l118_323_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_323 = _zz_when_ArraySlice_l118_323_1[5:0];
  assign _zz_when_ArraySlice_l173_323_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_323_1 = {1'd0, _zz_when_ArraySlice_l173_323_2};
  assign _zz_when_ArraySlice_l173_323_3 = (_zz_when_ArraySlice_l173_323_4 + _zz_when_ArraySlice_l173_323_9);
  assign _zz_when_ArraySlice_l173_323_4 = (_zz_when_ArraySlice_l173_323 - _zz_when_ArraySlice_l173_323_5);
  assign _zz_when_ArraySlice_l173_323_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_323_7);
  assign _zz_when_ArraySlice_l173_323_5 = {1'd0, _zz_when_ArraySlice_l173_323_6};
  assign _zz_when_ArraySlice_l173_323_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_323_7 = {1'd0, _zz_when_ArraySlice_l173_323_8};
  assign _zz_when_ArraySlice_l173_323_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_324 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_324_1);
  assign _zz_when_ArraySlice_l165_324_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_324 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_324_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_324_2);
  assign _zz_when_ArraySlice_l166_324_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_324_3);
  assign _zz_when_ArraySlice_l166_324_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_324 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_324 = (_zz_when_ArraySlice_l113_324_1 - _zz_when_ArraySlice_l113_324_4);
  assign _zz_when_ArraySlice_l113_324_1 = (_zz_when_ArraySlice_l113_324_2 + _zz_when_ArraySlice_l113_324_3);
  assign _zz_when_ArraySlice_l113_324_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_324_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_324_4 = {1'd0, _zz_when_ArraySlice_l112_324};
  assign _zz__zz_when_ArraySlice_l173_324 = (_zz__zz_when_ArraySlice_l173_324_1 + _zz__zz_when_ArraySlice_l173_324_2);
  assign _zz__zz_when_ArraySlice_l173_324_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_324_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_324_3 = {1'd0, _zz_when_ArraySlice_l112_324};
  assign _zz_when_ArraySlice_l118_324_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_324 = _zz_when_ArraySlice_l118_324_1[5:0];
  assign _zz_when_ArraySlice_l173_324_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_324_1 = {1'd0, _zz_when_ArraySlice_l173_324_2};
  assign _zz_when_ArraySlice_l173_324_3 = (_zz_when_ArraySlice_l173_324_4 + _zz_when_ArraySlice_l173_324_8);
  assign _zz_when_ArraySlice_l173_324_4 = (_zz_when_ArraySlice_l173_324 - _zz_when_ArraySlice_l173_324_5);
  assign _zz_when_ArraySlice_l173_324_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_324_7);
  assign _zz_when_ArraySlice_l173_324_5 = {1'd0, _zz_when_ArraySlice_l173_324_6};
  assign _zz_when_ArraySlice_l173_324_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_324_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_325 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_325_1);
  assign _zz_when_ArraySlice_l165_325_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_325_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_325 = {1'd0, _zz_when_ArraySlice_l166_325_1};
  assign _zz_when_ArraySlice_l166_325_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_325_3);
  assign _zz_when_ArraySlice_l166_325_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_325_4);
  assign _zz_when_ArraySlice_l166_325_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_325 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_325 = (_zz_when_ArraySlice_l113_325_1 - _zz_when_ArraySlice_l113_325_4);
  assign _zz_when_ArraySlice_l113_325_1 = (_zz_when_ArraySlice_l113_325_2 + _zz_when_ArraySlice_l113_325_3);
  assign _zz_when_ArraySlice_l113_325_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_325_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_325_4 = {1'd0, _zz_when_ArraySlice_l112_325};
  assign _zz__zz_when_ArraySlice_l173_325 = (_zz__zz_when_ArraySlice_l173_325_1 + _zz__zz_when_ArraySlice_l173_325_2);
  assign _zz__zz_when_ArraySlice_l173_325_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_325_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_325_3 = {1'd0, _zz_when_ArraySlice_l112_325};
  assign _zz_when_ArraySlice_l118_325_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_325 = _zz_when_ArraySlice_l118_325_1[5:0];
  assign _zz_when_ArraySlice_l173_325_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_325_1 = {2'd0, _zz_when_ArraySlice_l173_325_2};
  assign _zz_when_ArraySlice_l173_325_3 = (_zz_when_ArraySlice_l173_325_4 + _zz_when_ArraySlice_l173_325_8);
  assign _zz_when_ArraySlice_l173_325_4 = (_zz_when_ArraySlice_l173_325 - _zz_when_ArraySlice_l173_325_5);
  assign _zz_when_ArraySlice_l173_325_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_325_7);
  assign _zz_when_ArraySlice_l173_325_5 = {1'd0, _zz_when_ArraySlice_l173_325_6};
  assign _zz_when_ArraySlice_l173_325_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_325_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_326 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_326_1);
  assign _zz_when_ArraySlice_l165_326_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_326_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_326 = {1'd0, _zz_when_ArraySlice_l166_326_1};
  assign _zz_when_ArraySlice_l166_326_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_326_3);
  assign _zz_when_ArraySlice_l166_326_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_326_4);
  assign _zz_when_ArraySlice_l166_326_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_326 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_326 = (_zz_when_ArraySlice_l113_326_1 - _zz_when_ArraySlice_l113_326_4);
  assign _zz_when_ArraySlice_l113_326_1 = (_zz_when_ArraySlice_l113_326_2 + _zz_when_ArraySlice_l113_326_3);
  assign _zz_when_ArraySlice_l113_326_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_326_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_326_4 = {1'd0, _zz_when_ArraySlice_l112_326};
  assign _zz__zz_when_ArraySlice_l173_326 = (_zz__zz_when_ArraySlice_l173_326_1 + _zz__zz_when_ArraySlice_l173_326_2);
  assign _zz__zz_when_ArraySlice_l173_326_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_326_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_326_3 = {1'd0, _zz_when_ArraySlice_l112_326};
  assign _zz_when_ArraySlice_l118_326_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_326 = _zz_when_ArraySlice_l118_326_1[5:0];
  assign _zz_when_ArraySlice_l173_326_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_326_1 = {2'd0, _zz_when_ArraySlice_l173_326_2};
  assign _zz_when_ArraySlice_l173_326_3 = (_zz_when_ArraySlice_l173_326_4 + _zz_when_ArraySlice_l173_326_8);
  assign _zz_when_ArraySlice_l173_326_4 = (_zz_when_ArraySlice_l173_326 - _zz_when_ArraySlice_l173_326_5);
  assign _zz_when_ArraySlice_l173_326_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_326_7);
  assign _zz_when_ArraySlice_l173_326_5 = {1'd0, _zz_when_ArraySlice_l173_326_6};
  assign _zz_when_ArraySlice_l173_326_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_326_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_327 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_327_1);
  assign _zz_when_ArraySlice_l165_327_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_327_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_327 = {2'd0, _zz_when_ArraySlice_l166_327_1};
  assign _zz_when_ArraySlice_l166_327_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_327_3);
  assign _zz_when_ArraySlice_l166_327_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_327_4);
  assign _zz_when_ArraySlice_l166_327_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_327 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_327 = (_zz_when_ArraySlice_l113_327_1 - _zz_when_ArraySlice_l113_327_4);
  assign _zz_when_ArraySlice_l113_327_1 = (_zz_when_ArraySlice_l113_327_2 + _zz_when_ArraySlice_l113_327_3);
  assign _zz_when_ArraySlice_l113_327_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_327_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_327_4 = {1'd0, _zz_when_ArraySlice_l112_327};
  assign _zz__zz_when_ArraySlice_l173_327 = (_zz__zz_when_ArraySlice_l173_327_1 + _zz__zz_when_ArraySlice_l173_327_2);
  assign _zz__zz_when_ArraySlice_l173_327_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_327_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_327_3 = {1'd0, _zz_when_ArraySlice_l112_327};
  assign _zz_when_ArraySlice_l118_327_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_327 = _zz_when_ArraySlice_l118_327_1[5:0];
  assign _zz_when_ArraySlice_l173_327_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_327_1 = {3'd0, _zz_when_ArraySlice_l173_327_2};
  assign _zz_when_ArraySlice_l173_327_3 = (_zz_when_ArraySlice_l173_327_4 + _zz_when_ArraySlice_l173_327_8);
  assign _zz_when_ArraySlice_l173_327_4 = (_zz_when_ArraySlice_l173_327 - _zz_when_ArraySlice_l173_327_5);
  assign _zz_when_ArraySlice_l173_327_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_327_7);
  assign _zz_when_ArraySlice_l173_327_5 = {1'd0, _zz_when_ArraySlice_l173_327_6};
  assign _zz_when_ArraySlice_l173_327_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_327_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_4_63 = 1'b1;
  assign _zz_selectReadFifo_4_62 = {5'd0, _zz_selectReadFifo_4_63};
  assign _zz_when_ArraySlice_l315_4 = (_zz_when_ArraySlice_l315_4_1 % aReg);
  assign _zz_when_ArraySlice_l315_4_1 = (handshakeTimes_4_value + _zz_when_ArraySlice_l315_4_2);
  assign _zz_when_ArraySlice_l315_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l315_4_2 = {12'd0, _zz_when_ArraySlice_l315_4_3};
  assign _zz_when_ArraySlice_l301_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l301_4_1);
  assign _zz_when_ArraySlice_l301_4_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l322_4_2 = (_zz_when_ArraySlice_l322_4_3 - _zz_when_ArraySlice_l322_4_4);
  assign _zz_when_ArraySlice_l322_4_1 = {7'd0, _zz_when_ArraySlice_l322_4_2};
  assign _zz_when_ArraySlice_l322_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l322_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l322_4_4 = {5'd0, _zz_when_ArraySlice_l322_4_5};
  assign _zz_when_ArraySlice_l240_5 = (selectReadFifo_5 + _zz_when_ArraySlice_l240_5_1);
  assign _zz_when_ArraySlice_l240_5_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l241_5_1 = (selectReadFifo_5 + _zz_when_ArraySlice_l241_5_2);
  assign _zz_when_ArraySlice_l241_5_2 = (bReg * 3'b101);
  assign _zz__zz_outputStreamArrayData_5_valid_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l247_5_2 = 1'b1;
  assign _zz_when_ArraySlice_l247_5_1 = {6'd0, _zz_when_ArraySlice_l247_5_2};
  assign _zz_when_ArraySlice_l247_5_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l247_5_5);
  assign _zz_when_ArraySlice_l247_5_5 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l248_5_1 = (_zz_when_ArraySlice_l248_5_2 - _zz_when_ArraySlice_l248_5_3);
  assign _zz_when_ArraySlice_l248_5 = {7'd0, _zz_when_ArraySlice_l248_5_1};
  assign _zz_when_ArraySlice_l248_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l248_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l248_5_3 = {5'd0, _zz_when_ArraySlice_l248_5_4};
  assign _zz_selectReadFifo_5_32 = (selectReadFifo_5 - _zz_selectReadFifo_5_33);
  assign _zz_selectReadFifo_5_33 = {3'd0, bReg};
  assign _zz_selectReadFifo_5_35 = 1'b1;
  assign _zz_selectReadFifo_5_34 = {5'd0, _zz_selectReadFifo_5_35};
  assign _zz_selectReadFifo_5_37 = 1'b1;
  assign _zz_selectReadFifo_5_36 = {5'd0, _zz_selectReadFifo_5_37};
  assign _zz_when_ArraySlice_l251_5 = (_zz_when_ArraySlice_l251_5_1 % aReg);
  assign _zz_when_ArraySlice_l251_5_1 = (handshakeTimes_5_value + _zz_when_ArraySlice_l251_5_2);
  assign _zz_when_ArraySlice_l251_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l251_5_2 = {12'd0, _zz_when_ArraySlice_l251_5_3};
  assign _zz_when_ArraySlice_l256_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l256_5_3);
  assign _zz_when_ArraySlice_l256_5_3 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l256_5_5 = 1'b1;
  assign _zz_when_ArraySlice_l256_5_4 = {6'd0, _zz_when_ArraySlice_l256_5_5};
  assign _zz_when_ArraySlice_l257_5_1 = (_zz_when_ArraySlice_l257_5_2 - _zz_when_ArraySlice_l257_5_3);
  assign _zz_when_ArraySlice_l257_5 = {7'd0, _zz_when_ArraySlice_l257_5_1};
  assign _zz_when_ArraySlice_l257_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l257_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l257_5_3 = {5'd0, _zz_when_ArraySlice_l257_5_4};
  assign _zz__zz_when_ArraySlice_l94_39 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_39 = (_zz_when_ArraySlice_l95_39_1 - _zz_when_ArraySlice_l95_39_4);
  assign _zz_when_ArraySlice_l95_39_1 = (_zz_when_ArraySlice_l95_39_2 + _zz_when_ArraySlice_l95_39_3);
  assign _zz_when_ArraySlice_l95_39_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_39_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_39_4 = {1'd0, _zz_when_ArraySlice_l94_39};
  assign _zz__zz_when_ArraySlice_l259_5 = (_zz__zz_when_ArraySlice_l259_5_1 + _zz__zz_when_ArraySlice_l259_5_2);
  assign _zz__zz_when_ArraySlice_l259_5_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l259_5_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l259_5_3 = {1'd0, _zz_when_ArraySlice_l94_39};
  assign _zz_when_ArraySlice_l99_39_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_39 = _zz_when_ArraySlice_l99_39_1[5:0];
  assign _zz_when_ArraySlice_l259_5_1 = (outSliceNumb_5_value + _zz_when_ArraySlice_l259_5_2);
  assign _zz_when_ArraySlice_l259_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l259_5_2 = {6'd0, _zz_when_ArraySlice_l259_5_3};
  assign _zz_when_ArraySlice_l259_5_4 = (_zz_when_ArraySlice_l259_5 / aReg);
  assign _zz_selectReadFifo_5_38 = (selectReadFifo_5 - _zz_selectReadFifo_5_39);
  assign _zz_selectReadFifo_5_39 = {3'd0, bReg};
  assign _zz_selectReadFifo_5_41 = 1'b1;
  assign _zz_selectReadFifo_5_40 = {5'd0, _zz_selectReadFifo_5_41};
  assign _zz_selectReadFifo_5_42 = (selectReadFifo_5 + _zz_selectReadFifo_5_43);
  assign _zz_selectReadFifo_5_43 = (3'b111 * bReg);
  assign _zz_selectReadFifo_5_45 = 1'b1;
  assign _zz_selectReadFifo_5_44 = {5'd0, _zz_selectReadFifo_5_45};
  assign _zz_when_ArraySlice_l165_328 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_328_1);
  assign _zz_when_ArraySlice_l165_328_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_328_1 = {3'd0, _zz_when_ArraySlice_l165_328_2};
  assign _zz_when_ArraySlice_l166_328 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_328_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_328_3);
  assign _zz_when_ArraySlice_l166_328_1 = {1'd0, _zz_when_ArraySlice_l166_328_2};
  assign _zz_when_ArraySlice_l166_328_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_328_4);
  assign _zz_when_ArraySlice_l166_328_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_328_4 = {3'd0, _zz_when_ArraySlice_l166_328_5};
  assign _zz__zz_when_ArraySlice_l112_328 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_328 = (_zz_when_ArraySlice_l113_328_1 - _zz_when_ArraySlice_l113_328_4);
  assign _zz_when_ArraySlice_l113_328_1 = (_zz_when_ArraySlice_l113_328_2 + _zz_when_ArraySlice_l113_328_3);
  assign _zz_when_ArraySlice_l113_328_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_328_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_328_4 = {1'd0, _zz_when_ArraySlice_l112_328};
  assign _zz__zz_when_ArraySlice_l173_328 = (_zz__zz_when_ArraySlice_l173_328_1 + _zz__zz_when_ArraySlice_l173_328_2);
  assign _zz__zz_when_ArraySlice_l173_328_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_328_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_328_3 = {1'd0, _zz_when_ArraySlice_l112_328};
  assign _zz_when_ArraySlice_l118_328_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_328 = _zz_when_ArraySlice_l118_328_1[5:0];
  assign _zz_when_ArraySlice_l173_328_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_328_2 = (_zz_when_ArraySlice_l173_328_3 + _zz_when_ArraySlice_l173_328_8);
  assign _zz_when_ArraySlice_l173_328_3 = (_zz_when_ArraySlice_l173_328 - _zz_when_ArraySlice_l173_328_4);
  assign _zz_when_ArraySlice_l173_328_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_328_6);
  assign _zz_when_ArraySlice_l173_328_4 = {1'd0, _zz_when_ArraySlice_l173_328_5};
  assign _zz_when_ArraySlice_l173_328_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_328_6 = {3'd0, _zz_when_ArraySlice_l173_328_7};
  assign _zz_when_ArraySlice_l173_328_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_329 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_329_1);
  assign _zz_when_ArraySlice_l165_329_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_329_1 = {2'd0, _zz_when_ArraySlice_l165_329_2};
  assign _zz_when_ArraySlice_l166_329 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_329_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_329_2);
  assign _zz_when_ArraySlice_l166_329_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_329_3);
  assign _zz_when_ArraySlice_l166_329_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_329_3 = {2'd0, _zz_when_ArraySlice_l166_329_4};
  assign _zz__zz_when_ArraySlice_l112_329 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_329 = (_zz_when_ArraySlice_l113_329_1 - _zz_when_ArraySlice_l113_329_4);
  assign _zz_when_ArraySlice_l113_329_1 = (_zz_when_ArraySlice_l113_329_2 + _zz_when_ArraySlice_l113_329_3);
  assign _zz_when_ArraySlice_l113_329_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_329_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_329_4 = {1'd0, _zz_when_ArraySlice_l112_329};
  assign _zz__zz_when_ArraySlice_l173_329 = (_zz__zz_when_ArraySlice_l173_329_1 + _zz__zz_when_ArraySlice_l173_329_2);
  assign _zz__zz_when_ArraySlice_l173_329_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_329_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_329_3 = {1'd0, _zz_when_ArraySlice_l112_329};
  assign _zz_when_ArraySlice_l118_329_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_329 = _zz_when_ArraySlice_l118_329_1[5:0];
  assign _zz_when_ArraySlice_l173_329_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_329_1 = {1'd0, _zz_when_ArraySlice_l173_329_2};
  assign _zz_when_ArraySlice_l173_329_3 = (_zz_when_ArraySlice_l173_329_4 + _zz_when_ArraySlice_l173_329_9);
  assign _zz_when_ArraySlice_l173_329_4 = (_zz_when_ArraySlice_l173_329 - _zz_when_ArraySlice_l173_329_5);
  assign _zz_when_ArraySlice_l173_329_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_329_7);
  assign _zz_when_ArraySlice_l173_329_5 = {1'd0, _zz_when_ArraySlice_l173_329_6};
  assign _zz_when_ArraySlice_l173_329_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_329_7 = {2'd0, _zz_when_ArraySlice_l173_329_8};
  assign _zz_when_ArraySlice_l173_329_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_330 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_330_1);
  assign _zz_when_ArraySlice_l165_330_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_330_1 = {1'd0, _zz_when_ArraySlice_l165_330_2};
  assign _zz_when_ArraySlice_l166_330 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_330_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_330_2);
  assign _zz_when_ArraySlice_l166_330_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_330_3);
  assign _zz_when_ArraySlice_l166_330_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_330_3 = {1'd0, _zz_when_ArraySlice_l166_330_4};
  assign _zz__zz_when_ArraySlice_l112_330 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_330 = (_zz_when_ArraySlice_l113_330_1 - _zz_when_ArraySlice_l113_330_4);
  assign _zz_when_ArraySlice_l113_330_1 = (_zz_when_ArraySlice_l113_330_2 + _zz_when_ArraySlice_l113_330_3);
  assign _zz_when_ArraySlice_l113_330_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_330_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_330_4 = {1'd0, _zz_when_ArraySlice_l112_330};
  assign _zz__zz_when_ArraySlice_l173_330 = (_zz__zz_when_ArraySlice_l173_330_1 + _zz__zz_when_ArraySlice_l173_330_2);
  assign _zz__zz_when_ArraySlice_l173_330_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_330_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_330_3 = {1'd0, _zz_when_ArraySlice_l112_330};
  assign _zz_when_ArraySlice_l118_330_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_330 = _zz_when_ArraySlice_l118_330_1[5:0];
  assign _zz_when_ArraySlice_l173_330_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_330_1 = {1'd0, _zz_when_ArraySlice_l173_330_2};
  assign _zz_when_ArraySlice_l173_330_3 = (_zz_when_ArraySlice_l173_330_4 + _zz_when_ArraySlice_l173_330_9);
  assign _zz_when_ArraySlice_l173_330_4 = (_zz_when_ArraySlice_l173_330 - _zz_when_ArraySlice_l173_330_5);
  assign _zz_when_ArraySlice_l173_330_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_330_7);
  assign _zz_when_ArraySlice_l173_330_5 = {1'd0, _zz_when_ArraySlice_l173_330_6};
  assign _zz_when_ArraySlice_l173_330_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_330_7 = {1'd0, _zz_when_ArraySlice_l173_330_8};
  assign _zz_when_ArraySlice_l173_330_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_331 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_331_1);
  assign _zz_when_ArraySlice_l165_331_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_331_1 = {1'd0, _zz_when_ArraySlice_l165_331_2};
  assign _zz_when_ArraySlice_l166_331 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_331_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_331_2);
  assign _zz_when_ArraySlice_l166_331_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_331_3);
  assign _zz_when_ArraySlice_l166_331_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_331_3 = {1'd0, _zz_when_ArraySlice_l166_331_4};
  assign _zz__zz_when_ArraySlice_l112_331 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_331 = (_zz_when_ArraySlice_l113_331_1 - _zz_when_ArraySlice_l113_331_4);
  assign _zz_when_ArraySlice_l113_331_1 = (_zz_when_ArraySlice_l113_331_2 + _zz_when_ArraySlice_l113_331_3);
  assign _zz_when_ArraySlice_l113_331_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_331_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_331_4 = {1'd0, _zz_when_ArraySlice_l112_331};
  assign _zz__zz_when_ArraySlice_l173_331 = (_zz__zz_when_ArraySlice_l173_331_1 + _zz__zz_when_ArraySlice_l173_331_2);
  assign _zz__zz_when_ArraySlice_l173_331_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_331_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_331_3 = {1'd0, _zz_when_ArraySlice_l112_331};
  assign _zz_when_ArraySlice_l118_331_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_331 = _zz_when_ArraySlice_l118_331_1[5:0];
  assign _zz_when_ArraySlice_l173_331_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_331_1 = {1'd0, _zz_when_ArraySlice_l173_331_2};
  assign _zz_when_ArraySlice_l173_331_3 = (_zz_when_ArraySlice_l173_331_4 + _zz_when_ArraySlice_l173_331_9);
  assign _zz_when_ArraySlice_l173_331_4 = (_zz_when_ArraySlice_l173_331 - _zz_when_ArraySlice_l173_331_5);
  assign _zz_when_ArraySlice_l173_331_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_331_7);
  assign _zz_when_ArraySlice_l173_331_5 = {1'd0, _zz_when_ArraySlice_l173_331_6};
  assign _zz_when_ArraySlice_l173_331_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_331_7 = {1'd0, _zz_when_ArraySlice_l173_331_8};
  assign _zz_when_ArraySlice_l173_331_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_332 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_332_1);
  assign _zz_when_ArraySlice_l165_332_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_332 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_332_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_332_2);
  assign _zz_when_ArraySlice_l166_332_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_332_3);
  assign _zz_when_ArraySlice_l166_332_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_332 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_332 = (_zz_when_ArraySlice_l113_332_1 - _zz_when_ArraySlice_l113_332_4);
  assign _zz_when_ArraySlice_l113_332_1 = (_zz_when_ArraySlice_l113_332_2 + _zz_when_ArraySlice_l113_332_3);
  assign _zz_when_ArraySlice_l113_332_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_332_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_332_4 = {1'd0, _zz_when_ArraySlice_l112_332};
  assign _zz__zz_when_ArraySlice_l173_332 = (_zz__zz_when_ArraySlice_l173_332_1 + _zz__zz_when_ArraySlice_l173_332_2);
  assign _zz__zz_when_ArraySlice_l173_332_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_332_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_332_3 = {1'd0, _zz_when_ArraySlice_l112_332};
  assign _zz_when_ArraySlice_l118_332_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_332 = _zz_when_ArraySlice_l118_332_1[5:0];
  assign _zz_when_ArraySlice_l173_332_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_332_1 = {1'd0, _zz_when_ArraySlice_l173_332_2};
  assign _zz_when_ArraySlice_l173_332_3 = (_zz_when_ArraySlice_l173_332_4 + _zz_when_ArraySlice_l173_332_8);
  assign _zz_when_ArraySlice_l173_332_4 = (_zz_when_ArraySlice_l173_332 - _zz_when_ArraySlice_l173_332_5);
  assign _zz_when_ArraySlice_l173_332_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_332_7);
  assign _zz_when_ArraySlice_l173_332_5 = {1'd0, _zz_when_ArraySlice_l173_332_6};
  assign _zz_when_ArraySlice_l173_332_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_332_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_333 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_333_1);
  assign _zz_when_ArraySlice_l165_333_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_333_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_333 = {1'd0, _zz_when_ArraySlice_l166_333_1};
  assign _zz_when_ArraySlice_l166_333_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_333_3);
  assign _zz_when_ArraySlice_l166_333_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_333_4);
  assign _zz_when_ArraySlice_l166_333_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_333 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_333 = (_zz_when_ArraySlice_l113_333_1 - _zz_when_ArraySlice_l113_333_4);
  assign _zz_when_ArraySlice_l113_333_1 = (_zz_when_ArraySlice_l113_333_2 + _zz_when_ArraySlice_l113_333_3);
  assign _zz_when_ArraySlice_l113_333_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_333_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_333_4 = {1'd0, _zz_when_ArraySlice_l112_333};
  assign _zz__zz_when_ArraySlice_l173_333 = (_zz__zz_when_ArraySlice_l173_333_1 + _zz__zz_when_ArraySlice_l173_333_2);
  assign _zz__zz_when_ArraySlice_l173_333_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_333_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_333_3 = {1'd0, _zz_when_ArraySlice_l112_333};
  assign _zz_when_ArraySlice_l118_333_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_333 = _zz_when_ArraySlice_l118_333_1[5:0];
  assign _zz_when_ArraySlice_l173_333_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_333_1 = {2'd0, _zz_when_ArraySlice_l173_333_2};
  assign _zz_when_ArraySlice_l173_333_3 = (_zz_when_ArraySlice_l173_333_4 + _zz_when_ArraySlice_l173_333_8);
  assign _zz_when_ArraySlice_l173_333_4 = (_zz_when_ArraySlice_l173_333 - _zz_when_ArraySlice_l173_333_5);
  assign _zz_when_ArraySlice_l173_333_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_333_7);
  assign _zz_when_ArraySlice_l173_333_5 = {1'd0, _zz_when_ArraySlice_l173_333_6};
  assign _zz_when_ArraySlice_l173_333_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_333_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_334 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_334_1);
  assign _zz_when_ArraySlice_l165_334_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_334_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_334 = {1'd0, _zz_when_ArraySlice_l166_334_1};
  assign _zz_when_ArraySlice_l166_334_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_334_3);
  assign _zz_when_ArraySlice_l166_334_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_334_4);
  assign _zz_when_ArraySlice_l166_334_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_334 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_334 = (_zz_when_ArraySlice_l113_334_1 - _zz_when_ArraySlice_l113_334_4);
  assign _zz_when_ArraySlice_l113_334_1 = (_zz_when_ArraySlice_l113_334_2 + _zz_when_ArraySlice_l113_334_3);
  assign _zz_when_ArraySlice_l113_334_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_334_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_334_4 = {1'd0, _zz_when_ArraySlice_l112_334};
  assign _zz__zz_when_ArraySlice_l173_334 = (_zz__zz_when_ArraySlice_l173_334_1 + _zz__zz_when_ArraySlice_l173_334_2);
  assign _zz__zz_when_ArraySlice_l173_334_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_334_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_334_3 = {1'd0, _zz_when_ArraySlice_l112_334};
  assign _zz_when_ArraySlice_l118_334_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_334 = _zz_when_ArraySlice_l118_334_1[5:0];
  assign _zz_when_ArraySlice_l173_334_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_334_1 = {2'd0, _zz_when_ArraySlice_l173_334_2};
  assign _zz_when_ArraySlice_l173_334_3 = (_zz_when_ArraySlice_l173_334_4 + _zz_when_ArraySlice_l173_334_8);
  assign _zz_when_ArraySlice_l173_334_4 = (_zz_when_ArraySlice_l173_334 - _zz_when_ArraySlice_l173_334_5);
  assign _zz_when_ArraySlice_l173_334_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_334_7);
  assign _zz_when_ArraySlice_l173_334_5 = {1'd0, _zz_when_ArraySlice_l173_334_6};
  assign _zz_when_ArraySlice_l173_334_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_334_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_335 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_335_1);
  assign _zz_when_ArraySlice_l165_335_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_335_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_335 = {2'd0, _zz_when_ArraySlice_l166_335_1};
  assign _zz_when_ArraySlice_l166_335_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_335_3);
  assign _zz_when_ArraySlice_l166_335_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_335_4);
  assign _zz_when_ArraySlice_l166_335_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_335 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_335 = (_zz_when_ArraySlice_l113_335_1 - _zz_when_ArraySlice_l113_335_4);
  assign _zz_when_ArraySlice_l113_335_1 = (_zz_when_ArraySlice_l113_335_2 + _zz_when_ArraySlice_l113_335_3);
  assign _zz_when_ArraySlice_l113_335_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_335_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_335_4 = {1'd0, _zz_when_ArraySlice_l112_335};
  assign _zz__zz_when_ArraySlice_l173_335 = (_zz__zz_when_ArraySlice_l173_335_1 + _zz__zz_when_ArraySlice_l173_335_2);
  assign _zz__zz_when_ArraySlice_l173_335_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_335_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_335_3 = {1'd0, _zz_when_ArraySlice_l112_335};
  assign _zz_when_ArraySlice_l118_335_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_335 = _zz_when_ArraySlice_l118_335_1[5:0];
  assign _zz_when_ArraySlice_l173_335_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_335_1 = {3'd0, _zz_when_ArraySlice_l173_335_2};
  assign _zz_when_ArraySlice_l173_335_3 = (_zz_when_ArraySlice_l173_335_4 + _zz_when_ArraySlice_l173_335_8);
  assign _zz_when_ArraySlice_l173_335_4 = (_zz_when_ArraySlice_l173_335 - _zz_when_ArraySlice_l173_335_5);
  assign _zz_when_ArraySlice_l173_335_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_335_7);
  assign _zz_when_ArraySlice_l173_335_5 = {1'd0, _zz_when_ArraySlice_l173_335_6};
  assign _zz_when_ArraySlice_l173_335_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_335_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l268_5_1 = (_zz_when_ArraySlice_l268_5_2 + _zz_when_ArraySlice_l268_5_7);
  assign _zz_when_ArraySlice_l268_5_2 = (_zz_when_ArraySlice_l268_5_3 + _zz_when_ArraySlice_l268_5_5);
  assign _zz_when_ArraySlice_l268_5_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l268_5_4);
  assign _zz_when_ArraySlice_l268_5_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l268_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l268_5_5 = {5'd0, _zz_when_ArraySlice_l268_5_6};
  assign _zz_when_ArraySlice_l268_5_7 = (bReg * 3'b101);
  assign _zz_selectReadFifo_5_47 = 1'b1;
  assign _zz_selectReadFifo_5_46 = {5'd0, _zz_selectReadFifo_5_47};
  assign _zz_when_ArraySlice_l272_5 = (_zz_when_ArraySlice_l272_5_1 % aReg);
  assign _zz_when_ArraySlice_l272_5_1 = (handshakeTimes_5_value + _zz_when_ArraySlice_l272_5_2);
  assign _zz_when_ArraySlice_l272_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l272_5_2 = {12'd0, _zz_when_ArraySlice_l272_5_3};
  assign _zz_when_ArraySlice_l276_5_1 = (selectReadFifo_5 + _zz_when_ArraySlice_l276_5_2);
  assign _zz_when_ArraySlice_l276_5_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l277_5_1 = (_zz_when_ArraySlice_l277_5_2 - _zz_when_ArraySlice_l277_5_3);
  assign _zz_when_ArraySlice_l277_5 = {7'd0, _zz_when_ArraySlice_l277_5_1};
  assign _zz_when_ArraySlice_l277_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l277_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l277_5_3 = {5'd0, _zz_when_ArraySlice_l277_5_4};
  assign _zz__zz_when_ArraySlice_l94_40 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_40 = (_zz_when_ArraySlice_l95_40_1 - _zz_when_ArraySlice_l95_40_4);
  assign _zz_when_ArraySlice_l95_40_1 = (_zz_when_ArraySlice_l95_40_2 + _zz_when_ArraySlice_l95_40_3);
  assign _zz_when_ArraySlice_l95_40_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_40_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_40_4 = {1'd0, _zz_when_ArraySlice_l94_40};
  assign _zz__zz_when_ArraySlice_l279_5 = (_zz__zz_when_ArraySlice_l279_5_1 + _zz__zz_when_ArraySlice_l279_5_2);
  assign _zz__zz_when_ArraySlice_l279_5_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l279_5_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l279_5_3 = {1'd0, _zz_when_ArraySlice_l94_40};
  assign _zz_when_ArraySlice_l99_40_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_40 = _zz_when_ArraySlice_l99_40_1[5:0];
  assign _zz_when_ArraySlice_l279_5_1 = (outSliceNumb_5_value + _zz_when_ArraySlice_l279_5_2);
  assign _zz_when_ArraySlice_l279_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l279_5_2 = {6'd0, _zz_when_ArraySlice_l279_5_3};
  assign _zz_when_ArraySlice_l279_5_4 = (_zz_when_ArraySlice_l279_5 / aReg);
  assign _zz_selectReadFifo_5_48 = (selectReadFifo_5 - _zz_selectReadFifo_5_49);
  assign _zz_selectReadFifo_5_49 = {3'd0, bReg};
  assign _zz_selectReadFifo_5_51 = 1'b1;
  assign _zz_selectReadFifo_5_50 = {5'd0, _zz_selectReadFifo_5_51};
  assign _zz_selectReadFifo_5_52 = (selectReadFifo_5 + _zz_selectReadFifo_5_53);
  assign _zz_selectReadFifo_5_53 = (3'b111 * bReg);
  assign _zz_selectReadFifo_5_55 = 1'b1;
  assign _zz_selectReadFifo_5_54 = {5'd0, _zz_selectReadFifo_5_55};
  assign _zz_when_ArraySlice_l165_336 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_336_1);
  assign _zz_when_ArraySlice_l165_336_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_336_1 = {3'd0, _zz_when_ArraySlice_l165_336_2};
  assign _zz_when_ArraySlice_l166_336 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_336_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_336_3);
  assign _zz_when_ArraySlice_l166_336_1 = {1'd0, _zz_when_ArraySlice_l166_336_2};
  assign _zz_when_ArraySlice_l166_336_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_336_4);
  assign _zz_when_ArraySlice_l166_336_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_336_4 = {3'd0, _zz_when_ArraySlice_l166_336_5};
  assign _zz__zz_when_ArraySlice_l112_336 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_336 = (_zz_when_ArraySlice_l113_336_1 - _zz_when_ArraySlice_l113_336_4);
  assign _zz_when_ArraySlice_l113_336_1 = (_zz_when_ArraySlice_l113_336_2 + _zz_when_ArraySlice_l113_336_3);
  assign _zz_when_ArraySlice_l113_336_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_336_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_336_4 = {1'd0, _zz_when_ArraySlice_l112_336};
  assign _zz__zz_when_ArraySlice_l173_336 = (_zz__zz_when_ArraySlice_l173_336_1 + _zz__zz_when_ArraySlice_l173_336_2);
  assign _zz__zz_when_ArraySlice_l173_336_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_336_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_336_3 = {1'd0, _zz_when_ArraySlice_l112_336};
  assign _zz_when_ArraySlice_l118_336_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_336 = _zz_when_ArraySlice_l118_336_1[5:0];
  assign _zz_when_ArraySlice_l173_336_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_336_2 = (_zz_when_ArraySlice_l173_336_3 + _zz_when_ArraySlice_l173_336_8);
  assign _zz_when_ArraySlice_l173_336_3 = (_zz_when_ArraySlice_l173_336 - _zz_when_ArraySlice_l173_336_4);
  assign _zz_when_ArraySlice_l173_336_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_336_6);
  assign _zz_when_ArraySlice_l173_336_4 = {1'd0, _zz_when_ArraySlice_l173_336_5};
  assign _zz_when_ArraySlice_l173_336_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_336_6 = {3'd0, _zz_when_ArraySlice_l173_336_7};
  assign _zz_when_ArraySlice_l173_336_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_337 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_337_1);
  assign _zz_when_ArraySlice_l165_337_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_337_1 = {2'd0, _zz_when_ArraySlice_l165_337_2};
  assign _zz_when_ArraySlice_l166_337 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_337_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_337_2);
  assign _zz_when_ArraySlice_l166_337_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_337_3);
  assign _zz_when_ArraySlice_l166_337_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_337_3 = {2'd0, _zz_when_ArraySlice_l166_337_4};
  assign _zz__zz_when_ArraySlice_l112_337 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_337 = (_zz_when_ArraySlice_l113_337_1 - _zz_when_ArraySlice_l113_337_4);
  assign _zz_when_ArraySlice_l113_337_1 = (_zz_when_ArraySlice_l113_337_2 + _zz_when_ArraySlice_l113_337_3);
  assign _zz_when_ArraySlice_l113_337_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_337_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_337_4 = {1'd0, _zz_when_ArraySlice_l112_337};
  assign _zz__zz_when_ArraySlice_l173_337 = (_zz__zz_when_ArraySlice_l173_337_1 + _zz__zz_when_ArraySlice_l173_337_2);
  assign _zz__zz_when_ArraySlice_l173_337_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_337_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_337_3 = {1'd0, _zz_when_ArraySlice_l112_337};
  assign _zz_when_ArraySlice_l118_337_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_337 = _zz_when_ArraySlice_l118_337_1[5:0];
  assign _zz_when_ArraySlice_l173_337_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_337_1 = {1'd0, _zz_when_ArraySlice_l173_337_2};
  assign _zz_when_ArraySlice_l173_337_3 = (_zz_when_ArraySlice_l173_337_4 + _zz_when_ArraySlice_l173_337_9);
  assign _zz_when_ArraySlice_l173_337_4 = (_zz_when_ArraySlice_l173_337 - _zz_when_ArraySlice_l173_337_5);
  assign _zz_when_ArraySlice_l173_337_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_337_7);
  assign _zz_when_ArraySlice_l173_337_5 = {1'd0, _zz_when_ArraySlice_l173_337_6};
  assign _zz_when_ArraySlice_l173_337_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_337_7 = {2'd0, _zz_when_ArraySlice_l173_337_8};
  assign _zz_when_ArraySlice_l173_337_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_338 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_338_1);
  assign _zz_when_ArraySlice_l165_338_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_338_1 = {1'd0, _zz_when_ArraySlice_l165_338_2};
  assign _zz_when_ArraySlice_l166_338 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_338_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_338_2);
  assign _zz_when_ArraySlice_l166_338_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_338_3);
  assign _zz_when_ArraySlice_l166_338_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_338_3 = {1'd0, _zz_when_ArraySlice_l166_338_4};
  assign _zz__zz_when_ArraySlice_l112_338 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_338 = (_zz_when_ArraySlice_l113_338_1 - _zz_when_ArraySlice_l113_338_4);
  assign _zz_when_ArraySlice_l113_338_1 = (_zz_when_ArraySlice_l113_338_2 + _zz_when_ArraySlice_l113_338_3);
  assign _zz_when_ArraySlice_l113_338_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_338_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_338_4 = {1'd0, _zz_when_ArraySlice_l112_338};
  assign _zz__zz_when_ArraySlice_l173_338 = (_zz__zz_when_ArraySlice_l173_338_1 + _zz__zz_when_ArraySlice_l173_338_2);
  assign _zz__zz_when_ArraySlice_l173_338_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_338_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_338_3 = {1'd0, _zz_when_ArraySlice_l112_338};
  assign _zz_when_ArraySlice_l118_338_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_338 = _zz_when_ArraySlice_l118_338_1[5:0];
  assign _zz_when_ArraySlice_l173_338_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_338_1 = {1'd0, _zz_when_ArraySlice_l173_338_2};
  assign _zz_when_ArraySlice_l173_338_3 = (_zz_when_ArraySlice_l173_338_4 + _zz_when_ArraySlice_l173_338_9);
  assign _zz_when_ArraySlice_l173_338_4 = (_zz_when_ArraySlice_l173_338 - _zz_when_ArraySlice_l173_338_5);
  assign _zz_when_ArraySlice_l173_338_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_338_7);
  assign _zz_when_ArraySlice_l173_338_5 = {1'd0, _zz_when_ArraySlice_l173_338_6};
  assign _zz_when_ArraySlice_l173_338_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_338_7 = {1'd0, _zz_when_ArraySlice_l173_338_8};
  assign _zz_when_ArraySlice_l173_338_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_339 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_339_1);
  assign _zz_when_ArraySlice_l165_339_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_339_1 = {1'd0, _zz_when_ArraySlice_l165_339_2};
  assign _zz_when_ArraySlice_l166_339 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_339_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_339_2);
  assign _zz_when_ArraySlice_l166_339_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_339_3);
  assign _zz_when_ArraySlice_l166_339_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_339_3 = {1'd0, _zz_when_ArraySlice_l166_339_4};
  assign _zz__zz_when_ArraySlice_l112_339 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_339 = (_zz_when_ArraySlice_l113_339_1 - _zz_when_ArraySlice_l113_339_4);
  assign _zz_when_ArraySlice_l113_339_1 = (_zz_when_ArraySlice_l113_339_2 + _zz_when_ArraySlice_l113_339_3);
  assign _zz_when_ArraySlice_l113_339_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_339_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_339_4 = {1'd0, _zz_when_ArraySlice_l112_339};
  assign _zz__zz_when_ArraySlice_l173_339 = (_zz__zz_when_ArraySlice_l173_339_1 + _zz__zz_when_ArraySlice_l173_339_2);
  assign _zz__zz_when_ArraySlice_l173_339_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_339_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_339_3 = {1'd0, _zz_when_ArraySlice_l112_339};
  assign _zz_when_ArraySlice_l118_339_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_339 = _zz_when_ArraySlice_l118_339_1[5:0];
  assign _zz_when_ArraySlice_l173_339_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_339_1 = {1'd0, _zz_when_ArraySlice_l173_339_2};
  assign _zz_when_ArraySlice_l173_339_3 = (_zz_when_ArraySlice_l173_339_4 + _zz_when_ArraySlice_l173_339_9);
  assign _zz_when_ArraySlice_l173_339_4 = (_zz_when_ArraySlice_l173_339 - _zz_when_ArraySlice_l173_339_5);
  assign _zz_when_ArraySlice_l173_339_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_339_7);
  assign _zz_when_ArraySlice_l173_339_5 = {1'd0, _zz_when_ArraySlice_l173_339_6};
  assign _zz_when_ArraySlice_l173_339_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_339_7 = {1'd0, _zz_when_ArraySlice_l173_339_8};
  assign _zz_when_ArraySlice_l173_339_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_340 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_340_1);
  assign _zz_when_ArraySlice_l165_340_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_340 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_340_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_340_2);
  assign _zz_when_ArraySlice_l166_340_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_340_3);
  assign _zz_when_ArraySlice_l166_340_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_340 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_340 = (_zz_when_ArraySlice_l113_340_1 - _zz_when_ArraySlice_l113_340_4);
  assign _zz_when_ArraySlice_l113_340_1 = (_zz_when_ArraySlice_l113_340_2 + _zz_when_ArraySlice_l113_340_3);
  assign _zz_when_ArraySlice_l113_340_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_340_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_340_4 = {1'd0, _zz_when_ArraySlice_l112_340};
  assign _zz__zz_when_ArraySlice_l173_340 = (_zz__zz_when_ArraySlice_l173_340_1 + _zz__zz_when_ArraySlice_l173_340_2);
  assign _zz__zz_when_ArraySlice_l173_340_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_340_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_340_3 = {1'd0, _zz_when_ArraySlice_l112_340};
  assign _zz_when_ArraySlice_l118_340_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_340 = _zz_when_ArraySlice_l118_340_1[5:0];
  assign _zz_when_ArraySlice_l173_340_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_340_1 = {1'd0, _zz_when_ArraySlice_l173_340_2};
  assign _zz_when_ArraySlice_l173_340_3 = (_zz_when_ArraySlice_l173_340_4 + _zz_when_ArraySlice_l173_340_8);
  assign _zz_when_ArraySlice_l173_340_4 = (_zz_when_ArraySlice_l173_340 - _zz_when_ArraySlice_l173_340_5);
  assign _zz_when_ArraySlice_l173_340_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_340_7);
  assign _zz_when_ArraySlice_l173_340_5 = {1'd0, _zz_when_ArraySlice_l173_340_6};
  assign _zz_when_ArraySlice_l173_340_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_340_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_341 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_341_1);
  assign _zz_when_ArraySlice_l165_341_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_341_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_341 = {1'd0, _zz_when_ArraySlice_l166_341_1};
  assign _zz_when_ArraySlice_l166_341_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_341_3);
  assign _zz_when_ArraySlice_l166_341_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_341_4);
  assign _zz_when_ArraySlice_l166_341_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_341 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_341 = (_zz_when_ArraySlice_l113_341_1 - _zz_when_ArraySlice_l113_341_4);
  assign _zz_when_ArraySlice_l113_341_1 = (_zz_when_ArraySlice_l113_341_2 + _zz_when_ArraySlice_l113_341_3);
  assign _zz_when_ArraySlice_l113_341_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_341_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_341_4 = {1'd0, _zz_when_ArraySlice_l112_341};
  assign _zz__zz_when_ArraySlice_l173_341 = (_zz__zz_when_ArraySlice_l173_341_1 + _zz__zz_when_ArraySlice_l173_341_2);
  assign _zz__zz_when_ArraySlice_l173_341_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_341_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_341_3 = {1'd0, _zz_when_ArraySlice_l112_341};
  assign _zz_when_ArraySlice_l118_341_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_341 = _zz_when_ArraySlice_l118_341_1[5:0];
  assign _zz_when_ArraySlice_l173_341_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_341_1 = {2'd0, _zz_when_ArraySlice_l173_341_2};
  assign _zz_when_ArraySlice_l173_341_3 = (_zz_when_ArraySlice_l173_341_4 + _zz_when_ArraySlice_l173_341_8);
  assign _zz_when_ArraySlice_l173_341_4 = (_zz_when_ArraySlice_l173_341 - _zz_when_ArraySlice_l173_341_5);
  assign _zz_when_ArraySlice_l173_341_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_341_7);
  assign _zz_when_ArraySlice_l173_341_5 = {1'd0, _zz_when_ArraySlice_l173_341_6};
  assign _zz_when_ArraySlice_l173_341_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_341_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_342 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_342_1);
  assign _zz_when_ArraySlice_l165_342_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_342_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_342 = {1'd0, _zz_when_ArraySlice_l166_342_1};
  assign _zz_when_ArraySlice_l166_342_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_342_3);
  assign _zz_when_ArraySlice_l166_342_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_342_4);
  assign _zz_when_ArraySlice_l166_342_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_342 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_342 = (_zz_when_ArraySlice_l113_342_1 - _zz_when_ArraySlice_l113_342_4);
  assign _zz_when_ArraySlice_l113_342_1 = (_zz_when_ArraySlice_l113_342_2 + _zz_when_ArraySlice_l113_342_3);
  assign _zz_when_ArraySlice_l113_342_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_342_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_342_4 = {1'd0, _zz_when_ArraySlice_l112_342};
  assign _zz__zz_when_ArraySlice_l173_342 = (_zz__zz_when_ArraySlice_l173_342_1 + _zz__zz_when_ArraySlice_l173_342_2);
  assign _zz__zz_when_ArraySlice_l173_342_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_342_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_342_3 = {1'd0, _zz_when_ArraySlice_l112_342};
  assign _zz_when_ArraySlice_l118_342_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_342 = _zz_when_ArraySlice_l118_342_1[5:0];
  assign _zz_when_ArraySlice_l173_342_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_342_1 = {2'd0, _zz_when_ArraySlice_l173_342_2};
  assign _zz_when_ArraySlice_l173_342_3 = (_zz_when_ArraySlice_l173_342_4 + _zz_when_ArraySlice_l173_342_8);
  assign _zz_when_ArraySlice_l173_342_4 = (_zz_when_ArraySlice_l173_342 - _zz_when_ArraySlice_l173_342_5);
  assign _zz_when_ArraySlice_l173_342_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_342_7);
  assign _zz_when_ArraySlice_l173_342_5 = {1'd0, _zz_when_ArraySlice_l173_342_6};
  assign _zz_when_ArraySlice_l173_342_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_342_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_343 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_343_1);
  assign _zz_when_ArraySlice_l165_343_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_343_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_343 = {2'd0, _zz_when_ArraySlice_l166_343_1};
  assign _zz_when_ArraySlice_l166_343_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_343_3);
  assign _zz_when_ArraySlice_l166_343_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_343_4);
  assign _zz_when_ArraySlice_l166_343_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_343 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_343 = (_zz_when_ArraySlice_l113_343_1 - _zz_when_ArraySlice_l113_343_4);
  assign _zz_when_ArraySlice_l113_343_1 = (_zz_when_ArraySlice_l113_343_2 + _zz_when_ArraySlice_l113_343_3);
  assign _zz_when_ArraySlice_l113_343_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_343_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_343_4 = {1'd0, _zz_when_ArraySlice_l112_343};
  assign _zz__zz_when_ArraySlice_l173_343 = (_zz__zz_when_ArraySlice_l173_343_1 + _zz__zz_when_ArraySlice_l173_343_2);
  assign _zz__zz_when_ArraySlice_l173_343_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_343_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_343_3 = {1'd0, _zz_when_ArraySlice_l112_343};
  assign _zz_when_ArraySlice_l118_343_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_343 = _zz_when_ArraySlice_l118_343_1[5:0];
  assign _zz_when_ArraySlice_l173_343_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_343_1 = {3'd0, _zz_when_ArraySlice_l173_343_2};
  assign _zz_when_ArraySlice_l173_343_3 = (_zz_when_ArraySlice_l173_343_4 + _zz_when_ArraySlice_l173_343_8);
  assign _zz_when_ArraySlice_l173_343_4 = (_zz_when_ArraySlice_l173_343 - _zz_when_ArraySlice_l173_343_5);
  assign _zz_when_ArraySlice_l173_343_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_343_7);
  assign _zz_when_ArraySlice_l173_343_5 = {1'd0, _zz_when_ArraySlice_l173_343_6};
  assign _zz_when_ArraySlice_l173_343_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_343_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l288_5_1 = (_zz_when_ArraySlice_l288_5_2 + _zz_when_ArraySlice_l288_5_7);
  assign _zz_when_ArraySlice_l288_5_2 = (_zz_when_ArraySlice_l288_5_3 + _zz_when_ArraySlice_l288_5_5);
  assign _zz_when_ArraySlice_l288_5_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l288_5_4);
  assign _zz_when_ArraySlice_l288_5_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l288_5_5 = {5'd0, _zz_when_ArraySlice_l288_5_6};
  assign _zz_when_ArraySlice_l288_5_7 = (bReg * 3'b101);
  assign _zz_selectReadFifo_5_57 = 1'b1;
  assign _zz_selectReadFifo_5_56 = {5'd0, _zz_selectReadFifo_5_57};
  assign _zz_when_ArraySlice_l292_5 = (_zz_when_ArraySlice_l292_5_1 % aReg);
  assign _zz_when_ArraySlice_l292_5_1 = (handshakeTimes_5_value + _zz_when_ArraySlice_l292_5_2);
  assign _zz_when_ArraySlice_l292_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l292_5_2 = {12'd0, _zz_when_ArraySlice_l292_5_3};
  assign _zz_when_ArraySlice_l303_5_1 = (_zz_when_ArraySlice_l303_5_2 - _zz_when_ArraySlice_l303_5_3);
  assign _zz_when_ArraySlice_l303_5 = {7'd0, _zz_when_ArraySlice_l303_5_1};
  assign _zz_when_ArraySlice_l303_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l303_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l303_5_3 = {5'd0, _zz_when_ArraySlice_l303_5_4};
  assign _zz__zz_when_ArraySlice_l94_41 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_41 = (_zz_when_ArraySlice_l95_41_1 - _zz_when_ArraySlice_l95_41_4);
  assign _zz_when_ArraySlice_l95_41_1 = (_zz_when_ArraySlice_l95_41_2 + _zz_when_ArraySlice_l95_41_3);
  assign _zz_when_ArraySlice_l95_41_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_41_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_41_4 = {1'd0, _zz_when_ArraySlice_l94_41};
  assign _zz__zz_when_ArraySlice_l304_5 = (_zz__zz_when_ArraySlice_l304_5_1 + _zz__zz_when_ArraySlice_l304_5_2);
  assign _zz__zz_when_ArraySlice_l304_5_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l304_5_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l304_5_3 = {1'd0, _zz_when_ArraySlice_l94_41};
  assign _zz_when_ArraySlice_l99_41_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_41 = _zz_when_ArraySlice_l99_41_1[5:0];
  assign _zz_when_ArraySlice_l304_5_1 = (outSliceNumb_5_value + _zz_when_ArraySlice_l304_5_2);
  assign _zz_when_ArraySlice_l304_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l304_5_2 = {6'd0, _zz_when_ArraySlice_l304_5_3};
  assign _zz_when_ArraySlice_l304_5_4 = (_zz_when_ArraySlice_l304_5 / aReg);
  assign _zz_selectReadFifo_5_58 = (selectReadFifo_5 - _zz_selectReadFifo_5_59);
  assign _zz_selectReadFifo_5_59 = {3'd0, bReg};
  assign _zz_selectReadFifo_5_61 = 1'b1;
  assign _zz_selectReadFifo_5_60 = {5'd0, _zz_selectReadFifo_5_61};
  assign _zz_when_ArraySlice_l165_344 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_344_1);
  assign _zz_when_ArraySlice_l165_344_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_344_1 = {3'd0, _zz_when_ArraySlice_l165_344_2};
  assign _zz_when_ArraySlice_l166_344 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_344_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_344_3);
  assign _zz_when_ArraySlice_l166_344_1 = {1'd0, _zz_when_ArraySlice_l166_344_2};
  assign _zz_when_ArraySlice_l166_344_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_344_4);
  assign _zz_when_ArraySlice_l166_344_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_344_4 = {3'd0, _zz_when_ArraySlice_l166_344_5};
  assign _zz__zz_when_ArraySlice_l112_344 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_344 = (_zz_when_ArraySlice_l113_344_1 - _zz_when_ArraySlice_l113_344_4);
  assign _zz_when_ArraySlice_l113_344_1 = (_zz_when_ArraySlice_l113_344_2 + _zz_when_ArraySlice_l113_344_3);
  assign _zz_when_ArraySlice_l113_344_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_344_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_344_4 = {1'd0, _zz_when_ArraySlice_l112_344};
  assign _zz__zz_when_ArraySlice_l173_344 = (_zz__zz_when_ArraySlice_l173_344_1 + _zz__zz_when_ArraySlice_l173_344_2);
  assign _zz__zz_when_ArraySlice_l173_344_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_344_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_344_3 = {1'd0, _zz_when_ArraySlice_l112_344};
  assign _zz_when_ArraySlice_l118_344_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_344 = _zz_when_ArraySlice_l118_344_1[5:0];
  assign _zz_when_ArraySlice_l173_344_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_344_2 = (_zz_when_ArraySlice_l173_344_3 + _zz_when_ArraySlice_l173_344_8);
  assign _zz_when_ArraySlice_l173_344_3 = (_zz_when_ArraySlice_l173_344 - _zz_when_ArraySlice_l173_344_4);
  assign _zz_when_ArraySlice_l173_344_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_344_6);
  assign _zz_when_ArraySlice_l173_344_4 = {1'd0, _zz_when_ArraySlice_l173_344_5};
  assign _zz_when_ArraySlice_l173_344_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_344_6 = {3'd0, _zz_when_ArraySlice_l173_344_7};
  assign _zz_when_ArraySlice_l173_344_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_345 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_345_1);
  assign _zz_when_ArraySlice_l165_345_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_345_1 = {2'd0, _zz_when_ArraySlice_l165_345_2};
  assign _zz_when_ArraySlice_l166_345 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_345_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_345_2);
  assign _zz_when_ArraySlice_l166_345_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_345_3);
  assign _zz_when_ArraySlice_l166_345_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_345_3 = {2'd0, _zz_when_ArraySlice_l166_345_4};
  assign _zz__zz_when_ArraySlice_l112_345 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_345 = (_zz_when_ArraySlice_l113_345_1 - _zz_when_ArraySlice_l113_345_4);
  assign _zz_when_ArraySlice_l113_345_1 = (_zz_when_ArraySlice_l113_345_2 + _zz_when_ArraySlice_l113_345_3);
  assign _zz_when_ArraySlice_l113_345_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_345_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_345_4 = {1'd0, _zz_when_ArraySlice_l112_345};
  assign _zz__zz_when_ArraySlice_l173_345 = (_zz__zz_when_ArraySlice_l173_345_1 + _zz__zz_when_ArraySlice_l173_345_2);
  assign _zz__zz_when_ArraySlice_l173_345_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_345_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_345_3 = {1'd0, _zz_when_ArraySlice_l112_345};
  assign _zz_when_ArraySlice_l118_345_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_345 = _zz_when_ArraySlice_l118_345_1[5:0];
  assign _zz_when_ArraySlice_l173_345_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_345_1 = {1'd0, _zz_when_ArraySlice_l173_345_2};
  assign _zz_when_ArraySlice_l173_345_3 = (_zz_when_ArraySlice_l173_345_4 + _zz_when_ArraySlice_l173_345_9);
  assign _zz_when_ArraySlice_l173_345_4 = (_zz_when_ArraySlice_l173_345 - _zz_when_ArraySlice_l173_345_5);
  assign _zz_when_ArraySlice_l173_345_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_345_7);
  assign _zz_when_ArraySlice_l173_345_5 = {1'd0, _zz_when_ArraySlice_l173_345_6};
  assign _zz_when_ArraySlice_l173_345_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_345_7 = {2'd0, _zz_when_ArraySlice_l173_345_8};
  assign _zz_when_ArraySlice_l173_345_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_346 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_346_1);
  assign _zz_when_ArraySlice_l165_346_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_346_1 = {1'd0, _zz_when_ArraySlice_l165_346_2};
  assign _zz_when_ArraySlice_l166_346 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_346_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_346_2);
  assign _zz_when_ArraySlice_l166_346_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_346_3);
  assign _zz_when_ArraySlice_l166_346_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_346_3 = {1'd0, _zz_when_ArraySlice_l166_346_4};
  assign _zz__zz_when_ArraySlice_l112_346 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_346 = (_zz_when_ArraySlice_l113_346_1 - _zz_when_ArraySlice_l113_346_4);
  assign _zz_when_ArraySlice_l113_346_1 = (_zz_when_ArraySlice_l113_346_2 + _zz_when_ArraySlice_l113_346_3);
  assign _zz_when_ArraySlice_l113_346_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_346_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_346_4 = {1'd0, _zz_when_ArraySlice_l112_346};
  assign _zz__zz_when_ArraySlice_l173_346 = (_zz__zz_when_ArraySlice_l173_346_1 + _zz__zz_when_ArraySlice_l173_346_2);
  assign _zz__zz_when_ArraySlice_l173_346_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_346_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_346_3 = {1'd0, _zz_when_ArraySlice_l112_346};
  assign _zz_when_ArraySlice_l118_346_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_346 = _zz_when_ArraySlice_l118_346_1[5:0];
  assign _zz_when_ArraySlice_l173_346_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_346_1 = {1'd0, _zz_when_ArraySlice_l173_346_2};
  assign _zz_when_ArraySlice_l173_346_3 = (_zz_when_ArraySlice_l173_346_4 + _zz_when_ArraySlice_l173_346_9);
  assign _zz_when_ArraySlice_l173_346_4 = (_zz_when_ArraySlice_l173_346 - _zz_when_ArraySlice_l173_346_5);
  assign _zz_when_ArraySlice_l173_346_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_346_7);
  assign _zz_when_ArraySlice_l173_346_5 = {1'd0, _zz_when_ArraySlice_l173_346_6};
  assign _zz_when_ArraySlice_l173_346_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_346_7 = {1'd0, _zz_when_ArraySlice_l173_346_8};
  assign _zz_when_ArraySlice_l173_346_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_347 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_347_1);
  assign _zz_when_ArraySlice_l165_347_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_347_1 = {1'd0, _zz_when_ArraySlice_l165_347_2};
  assign _zz_when_ArraySlice_l166_347 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_347_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_347_2);
  assign _zz_when_ArraySlice_l166_347_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_347_3);
  assign _zz_when_ArraySlice_l166_347_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_347_3 = {1'd0, _zz_when_ArraySlice_l166_347_4};
  assign _zz__zz_when_ArraySlice_l112_347 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_347 = (_zz_when_ArraySlice_l113_347_1 - _zz_when_ArraySlice_l113_347_4);
  assign _zz_when_ArraySlice_l113_347_1 = (_zz_when_ArraySlice_l113_347_2 + _zz_when_ArraySlice_l113_347_3);
  assign _zz_when_ArraySlice_l113_347_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_347_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_347_4 = {1'd0, _zz_when_ArraySlice_l112_347};
  assign _zz__zz_when_ArraySlice_l173_347 = (_zz__zz_when_ArraySlice_l173_347_1 + _zz__zz_when_ArraySlice_l173_347_2);
  assign _zz__zz_when_ArraySlice_l173_347_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_347_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_347_3 = {1'd0, _zz_when_ArraySlice_l112_347};
  assign _zz_when_ArraySlice_l118_347_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_347 = _zz_when_ArraySlice_l118_347_1[5:0];
  assign _zz_when_ArraySlice_l173_347_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_347_1 = {1'd0, _zz_when_ArraySlice_l173_347_2};
  assign _zz_when_ArraySlice_l173_347_3 = (_zz_when_ArraySlice_l173_347_4 + _zz_when_ArraySlice_l173_347_9);
  assign _zz_when_ArraySlice_l173_347_4 = (_zz_when_ArraySlice_l173_347 - _zz_when_ArraySlice_l173_347_5);
  assign _zz_when_ArraySlice_l173_347_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_347_7);
  assign _zz_when_ArraySlice_l173_347_5 = {1'd0, _zz_when_ArraySlice_l173_347_6};
  assign _zz_when_ArraySlice_l173_347_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_347_7 = {1'd0, _zz_when_ArraySlice_l173_347_8};
  assign _zz_when_ArraySlice_l173_347_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_348 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_348_1);
  assign _zz_when_ArraySlice_l165_348_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_348 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_348_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_348_2);
  assign _zz_when_ArraySlice_l166_348_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_348_3);
  assign _zz_when_ArraySlice_l166_348_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_348 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_348 = (_zz_when_ArraySlice_l113_348_1 - _zz_when_ArraySlice_l113_348_4);
  assign _zz_when_ArraySlice_l113_348_1 = (_zz_when_ArraySlice_l113_348_2 + _zz_when_ArraySlice_l113_348_3);
  assign _zz_when_ArraySlice_l113_348_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_348_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_348_4 = {1'd0, _zz_when_ArraySlice_l112_348};
  assign _zz__zz_when_ArraySlice_l173_348 = (_zz__zz_when_ArraySlice_l173_348_1 + _zz__zz_when_ArraySlice_l173_348_2);
  assign _zz__zz_when_ArraySlice_l173_348_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_348_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_348_3 = {1'd0, _zz_when_ArraySlice_l112_348};
  assign _zz_when_ArraySlice_l118_348_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_348 = _zz_when_ArraySlice_l118_348_1[5:0];
  assign _zz_when_ArraySlice_l173_348_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_348_1 = {1'd0, _zz_when_ArraySlice_l173_348_2};
  assign _zz_when_ArraySlice_l173_348_3 = (_zz_when_ArraySlice_l173_348_4 + _zz_when_ArraySlice_l173_348_8);
  assign _zz_when_ArraySlice_l173_348_4 = (_zz_when_ArraySlice_l173_348 - _zz_when_ArraySlice_l173_348_5);
  assign _zz_when_ArraySlice_l173_348_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_348_7);
  assign _zz_when_ArraySlice_l173_348_5 = {1'd0, _zz_when_ArraySlice_l173_348_6};
  assign _zz_when_ArraySlice_l173_348_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_348_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_349 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_349_1);
  assign _zz_when_ArraySlice_l165_349_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_349_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_349 = {1'd0, _zz_when_ArraySlice_l166_349_1};
  assign _zz_when_ArraySlice_l166_349_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_349_3);
  assign _zz_when_ArraySlice_l166_349_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_349_4);
  assign _zz_when_ArraySlice_l166_349_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_349 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_349 = (_zz_when_ArraySlice_l113_349_1 - _zz_when_ArraySlice_l113_349_4);
  assign _zz_when_ArraySlice_l113_349_1 = (_zz_when_ArraySlice_l113_349_2 + _zz_when_ArraySlice_l113_349_3);
  assign _zz_when_ArraySlice_l113_349_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_349_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_349_4 = {1'd0, _zz_when_ArraySlice_l112_349};
  assign _zz__zz_when_ArraySlice_l173_349 = (_zz__zz_when_ArraySlice_l173_349_1 + _zz__zz_when_ArraySlice_l173_349_2);
  assign _zz__zz_when_ArraySlice_l173_349_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_349_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_349_3 = {1'd0, _zz_when_ArraySlice_l112_349};
  assign _zz_when_ArraySlice_l118_349_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_349 = _zz_when_ArraySlice_l118_349_1[5:0];
  assign _zz_when_ArraySlice_l173_349_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_349_1 = {2'd0, _zz_when_ArraySlice_l173_349_2};
  assign _zz_when_ArraySlice_l173_349_3 = (_zz_when_ArraySlice_l173_349_4 + _zz_when_ArraySlice_l173_349_8);
  assign _zz_when_ArraySlice_l173_349_4 = (_zz_when_ArraySlice_l173_349 - _zz_when_ArraySlice_l173_349_5);
  assign _zz_when_ArraySlice_l173_349_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_349_7);
  assign _zz_when_ArraySlice_l173_349_5 = {1'd0, _zz_when_ArraySlice_l173_349_6};
  assign _zz_when_ArraySlice_l173_349_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_349_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_350 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_350_1);
  assign _zz_when_ArraySlice_l165_350_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_350_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_350 = {1'd0, _zz_when_ArraySlice_l166_350_1};
  assign _zz_when_ArraySlice_l166_350_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_350_3);
  assign _zz_when_ArraySlice_l166_350_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_350_4);
  assign _zz_when_ArraySlice_l166_350_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_350 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_350 = (_zz_when_ArraySlice_l113_350_1 - _zz_when_ArraySlice_l113_350_4);
  assign _zz_when_ArraySlice_l113_350_1 = (_zz_when_ArraySlice_l113_350_2 + _zz_when_ArraySlice_l113_350_3);
  assign _zz_when_ArraySlice_l113_350_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_350_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_350_4 = {1'd0, _zz_when_ArraySlice_l112_350};
  assign _zz__zz_when_ArraySlice_l173_350 = (_zz__zz_when_ArraySlice_l173_350_1 + _zz__zz_when_ArraySlice_l173_350_2);
  assign _zz__zz_when_ArraySlice_l173_350_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_350_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_350_3 = {1'd0, _zz_when_ArraySlice_l112_350};
  assign _zz_when_ArraySlice_l118_350_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_350 = _zz_when_ArraySlice_l118_350_1[5:0];
  assign _zz_when_ArraySlice_l173_350_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_350_1 = {2'd0, _zz_when_ArraySlice_l173_350_2};
  assign _zz_when_ArraySlice_l173_350_3 = (_zz_when_ArraySlice_l173_350_4 + _zz_when_ArraySlice_l173_350_8);
  assign _zz_when_ArraySlice_l173_350_4 = (_zz_when_ArraySlice_l173_350 - _zz_when_ArraySlice_l173_350_5);
  assign _zz_when_ArraySlice_l173_350_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_350_7);
  assign _zz_when_ArraySlice_l173_350_5 = {1'd0, _zz_when_ArraySlice_l173_350_6};
  assign _zz_when_ArraySlice_l173_350_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_350_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_351 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_351_1);
  assign _zz_when_ArraySlice_l165_351_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_351_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_351 = {2'd0, _zz_when_ArraySlice_l166_351_1};
  assign _zz_when_ArraySlice_l166_351_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_351_3);
  assign _zz_when_ArraySlice_l166_351_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_351_4);
  assign _zz_when_ArraySlice_l166_351_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_351 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_351 = (_zz_when_ArraySlice_l113_351_1 - _zz_when_ArraySlice_l113_351_4);
  assign _zz_when_ArraySlice_l113_351_1 = (_zz_when_ArraySlice_l113_351_2 + _zz_when_ArraySlice_l113_351_3);
  assign _zz_when_ArraySlice_l113_351_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_351_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_351_4 = {1'd0, _zz_when_ArraySlice_l112_351};
  assign _zz__zz_when_ArraySlice_l173_351 = (_zz__zz_when_ArraySlice_l173_351_1 + _zz__zz_when_ArraySlice_l173_351_2);
  assign _zz__zz_when_ArraySlice_l173_351_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_351_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_351_3 = {1'd0, _zz_when_ArraySlice_l112_351};
  assign _zz_when_ArraySlice_l118_351_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_351 = _zz_when_ArraySlice_l118_351_1[5:0];
  assign _zz_when_ArraySlice_l173_351_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_351_1 = {3'd0, _zz_when_ArraySlice_l173_351_2};
  assign _zz_when_ArraySlice_l173_351_3 = (_zz_when_ArraySlice_l173_351_4 + _zz_when_ArraySlice_l173_351_8);
  assign _zz_when_ArraySlice_l173_351_4 = (_zz_when_ArraySlice_l173_351 - _zz_when_ArraySlice_l173_351_5);
  assign _zz_when_ArraySlice_l173_351_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_351_7);
  assign _zz_when_ArraySlice_l173_351_5 = {1'd0, _zz_when_ArraySlice_l173_351_6};
  assign _zz_when_ArraySlice_l173_351_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_351_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_5_63 = 1'b1;
  assign _zz_selectReadFifo_5_62 = {5'd0, _zz_selectReadFifo_5_63};
  assign _zz_when_ArraySlice_l315_5 = (_zz_when_ArraySlice_l315_5_1 % aReg);
  assign _zz_when_ArraySlice_l315_5_1 = (handshakeTimes_5_value + _zz_when_ArraySlice_l315_5_2);
  assign _zz_when_ArraySlice_l315_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l315_5_2 = {12'd0, _zz_when_ArraySlice_l315_5_3};
  assign _zz_when_ArraySlice_l301_5 = (selectReadFifo_5 + _zz_when_ArraySlice_l301_5_1);
  assign _zz_when_ArraySlice_l301_5_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l322_5_1 = (_zz_when_ArraySlice_l322_5_2 - _zz_when_ArraySlice_l322_5_3);
  assign _zz_when_ArraySlice_l322_5 = {7'd0, _zz_when_ArraySlice_l322_5_1};
  assign _zz_when_ArraySlice_l322_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l322_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l322_5_3 = {5'd0, _zz_when_ArraySlice_l322_5_4};
  assign _zz_when_ArraySlice_l240_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l240_6_1);
  assign _zz_when_ArraySlice_l240_6_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l241_6_1 = (selectReadFifo_6 + _zz_when_ArraySlice_l241_6_2);
  assign _zz_when_ArraySlice_l241_6_2 = (bReg * 3'b110);
  assign _zz__zz_outputStreamArrayData_6_valid_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l247_6_1 = 1'b1;
  assign _zz_when_ArraySlice_l247_6 = {6'd0, _zz_when_ArraySlice_l247_6_1};
  assign _zz_when_ArraySlice_l247_6_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l247_6_4);
  assign _zz_when_ArraySlice_l247_6_4 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l248_6_1 = (_zz_when_ArraySlice_l248_6_2 - _zz_when_ArraySlice_l248_6_3);
  assign _zz_when_ArraySlice_l248_6 = {7'd0, _zz_when_ArraySlice_l248_6_1};
  assign _zz_when_ArraySlice_l248_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l248_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l248_6_3 = {5'd0, _zz_when_ArraySlice_l248_6_4};
  assign _zz_selectReadFifo_6_32 = (selectReadFifo_6 - _zz_selectReadFifo_6_33);
  assign _zz_selectReadFifo_6_33 = {3'd0, bReg};
  assign _zz_selectReadFifo_6_35 = 1'b1;
  assign _zz_selectReadFifo_6_34 = {5'd0, _zz_selectReadFifo_6_35};
  assign _zz_selectReadFifo_6_37 = 1'b1;
  assign _zz_selectReadFifo_6_36 = {5'd0, _zz_selectReadFifo_6_37};
  assign _zz_when_ArraySlice_l251_6 = (_zz_when_ArraySlice_l251_6_1 % aReg);
  assign _zz_when_ArraySlice_l251_6_1 = (handshakeTimes_6_value + _zz_when_ArraySlice_l251_6_2);
  assign _zz_when_ArraySlice_l251_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l251_6_2 = {12'd0, _zz_when_ArraySlice_l251_6_3};
  assign _zz_when_ArraySlice_l256_6_1 = (selectReadFifo_6 + _zz_when_ArraySlice_l256_6_2);
  assign _zz_when_ArraySlice_l256_6_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l256_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l256_6_3 = {6'd0, _zz_when_ArraySlice_l256_6_4};
  assign _zz_when_ArraySlice_l257_6_1 = (_zz_when_ArraySlice_l257_6_2 - _zz_when_ArraySlice_l257_6_3);
  assign _zz_when_ArraySlice_l257_6 = {7'd0, _zz_when_ArraySlice_l257_6_1};
  assign _zz_when_ArraySlice_l257_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l257_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l257_6_3 = {5'd0, _zz_when_ArraySlice_l257_6_4};
  assign _zz__zz_when_ArraySlice_l94_42 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_42 = (_zz_when_ArraySlice_l95_42_1 - _zz_when_ArraySlice_l95_42_4);
  assign _zz_when_ArraySlice_l95_42_1 = (_zz_when_ArraySlice_l95_42_2 + _zz_when_ArraySlice_l95_42_3);
  assign _zz_when_ArraySlice_l95_42_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_42_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_42_4 = {1'd0, _zz_when_ArraySlice_l94_42};
  assign _zz__zz_when_ArraySlice_l259_6 = (_zz__zz_when_ArraySlice_l259_6_1 + _zz__zz_when_ArraySlice_l259_6_2);
  assign _zz__zz_when_ArraySlice_l259_6_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l259_6_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l259_6_3 = {1'd0, _zz_when_ArraySlice_l94_42};
  assign _zz_when_ArraySlice_l99_42_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_42 = _zz_when_ArraySlice_l99_42_1[5:0];
  assign _zz_when_ArraySlice_l259_6_1 = (outSliceNumb_6_value + _zz_when_ArraySlice_l259_6_2);
  assign _zz_when_ArraySlice_l259_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l259_6_2 = {6'd0, _zz_when_ArraySlice_l259_6_3};
  assign _zz_when_ArraySlice_l259_6_4 = (_zz_when_ArraySlice_l259_6 / aReg);
  assign _zz_selectReadFifo_6_38 = (selectReadFifo_6 - _zz_selectReadFifo_6_39);
  assign _zz_selectReadFifo_6_39 = {3'd0, bReg};
  assign _zz_selectReadFifo_6_41 = 1'b1;
  assign _zz_selectReadFifo_6_40 = {5'd0, _zz_selectReadFifo_6_41};
  assign _zz_selectReadFifo_6_42 = (selectReadFifo_6 + _zz_selectReadFifo_6_43);
  assign _zz_selectReadFifo_6_43 = (3'b111 * bReg);
  assign _zz_selectReadFifo_6_45 = 1'b1;
  assign _zz_selectReadFifo_6_44 = {5'd0, _zz_selectReadFifo_6_45};
  assign _zz_when_ArraySlice_l165_352 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_352_1);
  assign _zz_when_ArraySlice_l165_352_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_352_1 = {3'd0, _zz_when_ArraySlice_l165_352_2};
  assign _zz_when_ArraySlice_l166_352 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_352_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_352_3);
  assign _zz_when_ArraySlice_l166_352_1 = {1'd0, _zz_when_ArraySlice_l166_352_2};
  assign _zz_when_ArraySlice_l166_352_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_352_4);
  assign _zz_when_ArraySlice_l166_352_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_352_4 = {3'd0, _zz_when_ArraySlice_l166_352_5};
  assign _zz__zz_when_ArraySlice_l112_352 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_352 = (_zz_when_ArraySlice_l113_352_1 - _zz_when_ArraySlice_l113_352_4);
  assign _zz_when_ArraySlice_l113_352_1 = (_zz_when_ArraySlice_l113_352_2 + _zz_when_ArraySlice_l113_352_3);
  assign _zz_when_ArraySlice_l113_352_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_352_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_352_4 = {1'd0, _zz_when_ArraySlice_l112_352};
  assign _zz__zz_when_ArraySlice_l173_352 = (_zz__zz_when_ArraySlice_l173_352_1 + _zz__zz_when_ArraySlice_l173_352_2);
  assign _zz__zz_when_ArraySlice_l173_352_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_352_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_352_3 = {1'd0, _zz_when_ArraySlice_l112_352};
  assign _zz_when_ArraySlice_l118_352_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_352 = _zz_when_ArraySlice_l118_352_1[5:0];
  assign _zz_when_ArraySlice_l173_352_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_352_2 = (_zz_when_ArraySlice_l173_352_3 + _zz_when_ArraySlice_l173_352_8);
  assign _zz_when_ArraySlice_l173_352_3 = (_zz_when_ArraySlice_l173_352 - _zz_when_ArraySlice_l173_352_4);
  assign _zz_when_ArraySlice_l173_352_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_352_6);
  assign _zz_when_ArraySlice_l173_352_4 = {1'd0, _zz_when_ArraySlice_l173_352_5};
  assign _zz_when_ArraySlice_l173_352_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_352_6 = {3'd0, _zz_when_ArraySlice_l173_352_7};
  assign _zz_when_ArraySlice_l173_352_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_353 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_353_1);
  assign _zz_when_ArraySlice_l165_353_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_353_1 = {2'd0, _zz_when_ArraySlice_l165_353_2};
  assign _zz_when_ArraySlice_l166_353 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_353_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_353_2);
  assign _zz_when_ArraySlice_l166_353_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_353_3);
  assign _zz_when_ArraySlice_l166_353_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_353_3 = {2'd0, _zz_when_ArraySlice_l166_353_4};
  assign _zz__zz_when_ArraySlice_l112_353 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_353 = (_zz_when_ArraySlice_l113_353_1 - _zz_when_ArraySlice_l113_353_4);
  assign _zz_when_ArraySlice_l113_353_1 = (_zz_when_ArraySlice_l113_353_2 + _zz_when_ArraySlice_l113_353_3);
  assign _zz_when_ArraySlice_l113_353_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_353_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_353_4 = {1'd0, _zz_when_ArraySlice_l112_353};
  assign _zz__zz_when_ArraySlice_l173_353 = (_zz__zz_when_ArraySlice_l173_353_1 + _zz__zz_when_ArraySlice_l173_353_2);
  assign _zz__zz_when_ArraySlice_l173_353_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_353_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_353_3 = {1'd0, _zz_when_ArraySlice_l112_353};
  assign _zz_when_ArraySlice_l118_353_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_353 = _zz_when_ArraySlice_l118_353_1[5:0];
  assign _zz_when_ArraySlice_l173_353_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_353_1 = {1'd0, _zz_when_ArraySlice_l173_353_2};
  assign _zz_when_ArraySlice_l173_353_3 = (_zz_when_ArraySlice_l173_353_4 + _zz_when_ArraySlice_l173_353_9);
  assign _zz_when_ArraySlice_l173_353_4 = (_zz_when_ArraySlice_l173_353 - _zz_when_ArraySlice_l173_353_5);
  assign _zz_when_ArraySlice_l173_353_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_353_7);
  assign _zz_when_ArraySlice_l173_353_5 = {1'd0, _zz_when_ArraySlice_l173_353_6};
  assign _zz_when_ArraySlice_l173_353_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_353_7 = {2'd0, _zz_when_ArraySlice_l173_353_8};
  assign _zz_when_ArraySlice_l173_353_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_354 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_354_1);
  assign _zz_when_ArraySlice_l165_354_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_354_1 = {1'd0, _zz_when_ArraySlice_l165_354_2};
  assign _zz_when_ArraySlice_l166_354 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_354_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_354_2);
  assign _zz_when_ArraySlice_l166_354_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_354_3);
  assign _zz_when_ArraySlice_l166_354_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_354_3 = {1'd0, _zz_when_ArraySlice_l166_354_4};
  assign _zz__zz_when_ArraySlice_l112_354 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_354 = (_zz_when_ArraySlice_l113_354_1 - _zz_when_ArraySlice_l113_354_4);
  assign _zz_when_ArraySlice_l113_354_1 = (_zz_when_ArraySlice_l113_354_2 + _zz_when_ArraySlice_l113_354_3);
  assign _zz_when_ArraySlice_l113_354_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_354_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_354_4 = {1'd0, _zz_when_ArraySlice_l112_354};
  assign _zz__zz_when_ArraySlice_l173_354 = (_zz__zz_when_ArraySlice_l173_354_1 + _zz__zz_when_ArraySlice_l173_354_2);
  assign _zz__zz_when_ArraySlice_l173_354_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_354_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_354_3 = {1'd0, _zz_when_ArraySlice_l112_354};
  assign _zz_when_ArraySlice_l118_354_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_354 = _zz_when_ArraySlice_l118_354_1[5:0];
  assign _zz_when_ArraySlice_l173_354_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_354_1 = {1'd0, _zz_when_ArraySlice_l173_354_2};
  assign _zz_when_ArraySlice_l173_354_3 = (_zz_when_ArraySlice_l173_354_4 + _zz_when_ArraySlice_l173_354_9);
  assign _zz_when_ArraySlice_l173_354_4 = (_zz_when_ArraySlice_l173_354 - _zz_when_ArraySlice_l173_354_5);
  assign _zz_when_ArraySlice_l173_354_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_354_7);
  assign _zz_when_ArraySlice_l173_354_5 = {1'd0, _zz_when_ArraySlice_l173_354_6};
  assign _zz_when_ArraySlice_l173_354_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_354_7 = {1'd0, _zz_when_ArraySlice_l173_354_8};
  assign _zz_when_ArraySlice_l173_354_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_355 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_355_1);
  assign _zz_when_ArraySlice_l165_355_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_355_1 = {1'd0, _zz_when_ArraySlice_l165_355_2};
  assign _zz_when_ArraySlice_l166_355 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_355_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_355_2);
  assign _zz_when_ArraySlice_l166_355_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_355_3);
  assign _zz_when_ArraySlice_l166_355_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_355_3 = {1'd0, _zz_when_ArraySlice_l166_355_4};
  assign _zz__zz_when_ArraySlice_l112_355 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_355 = (_zz_when_ArraySlice_l113_355_1 - _zz_when_ArraySlice_l113_355_4);
  assign _zz_when_ArraySlice_l113_355_1 = (_zz_when_ArraySlice_l113_355_2 + _zz_when_ArraySlice_l113_355_3);
  assign _zz_when_ArraySlice_l113_355_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_355_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_355_4 = {1'd0, _zz_when_ArraySlice_l112_355};
  assign _zz__zz_when_ArraySlice_l173_355 = (_zz__zz_when_ArraySlice_l173_355_1 + _zz__zz_when_ArraySlice_l173_355_2);
  assign _zz__zz_when_ArraySlice_l173_355_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_355_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_355_3 = {1'd0, _zz_when_ArraySlice_l112_355};
  assign _zz_when_ArraySlice_l118_355_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_355 = _zz_when_ArraySlice_l118_355_1[5:0];
  assign _zz_when_ArraySlice_l173_355_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_355_1 = {1'd0, _zz_when_ArraySlice_l173_355_2};
  assign _zz_when_ArraySlice_l173_355_3 = (_zz_when_ArraySlice_l173_355_4 + _zz_when_ArraySlice_l173_355_9);
  assign _zz_when_ArraySlice_l173_355_4 = (_zz_when_ArraySlice_l173_355 - _zz_when_ArraySlice_l173_355_5);
  assign _zz_when_ArraySlice_l173_355_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_355_7);
  assign _zz_when_ArraySlice_l173_355_5 = {1'd0, _zz_when_ArraySlice_l173_355_6};
  assign _zz_when_ArraySlice_l173_355_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_355_7 = {1'd0, _zz_when_ArraySlice_l173_355_8};
  assign _zz_when_ArraySlice_l173_355_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_356 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_356_1);
  assign _zz_when_ArraySlice_l165_356_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_356 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_356_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_356_2);
  assign _zz_when_ArraySlice_l166_356_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_356_3);
  assign _zz_when_ArraySlice_l166_356_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_356 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_356 = (_zz_when_ArraySlice_l113_356_1 - _zz_when_ArraySlice_l113_356_4);
  assign _zz_when_ArraySlice_l113_356_1 = (_zz_when_ArraySlice_l113_356_2 + _zz_when_ArraySlice_l113_356_3);
  assign _zz_when_ArraySlice_l113_356_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_356_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_356_4 = {1'd0, _zz_when_ArraySlice_l112_356};
  assign _zz__zz_when_ArraySlice_l173_356 = (_zz__zz_when_ArraySlice_l173_356_1 + _zz__zz_when_ArraySlice_l173_356_2);
  assign _zz__zz_when_ArraySlice_l173_356_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_356_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_356_3 = {1'd0, _zz_when_ArraySlice_l112_356};
  assign _zz_when_ArraySlice_l118_356_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_356 = _zz_when_ArraySlice_l118_356_1[5:0];
  assign _zz_when_ArraySlice_l173_356_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_356_1 = {1'd0, _zz_when_ArraySlice_l173_356_2};
  assign _zz_when_ArraySlice_l173_356_3 = (_zz_when_ArraySlice_l173_356_4 + _zz_when_ArraySlice_l173_356_8);
  assign _zz_when_ArraySlice_l173_356_4 = (_zz_when_ArraySlice_l173_356 - _zz_when_ArraySlice_l173_356_5);
  assign _zz_when_ArraySlice_l173_356_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_356_7);
  assign _zz_when_ArraySlice_l173_356_5 = {1'd0, _zz_when_ArraySlice_l173_356_6};
  assign _zz_when_ArraySlice_l173_356_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_356_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_357 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_357_1);
  assign _zz_when_ArraySlice_l165_357_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_357_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_357 = {1'd0, _zz_when_ArraySlice_l166_357_1};
  assign _zz_when_ArraySlice_l166_357_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_357_3);
  assign _zz_when_ArraySlice_l166_357_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_357_4);
  assign _zz_when_ArraySlice_l166_357_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_357 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_357 = (_zz_when_ArraySlice_l113_357_1 - _zz_when_ArraySlice_l113_357_4);
  assign _zz_when_ArraySlice_l113_357_1 = (_zz_when_ArraySlice_l113_357_2 + _zz_when_ArraySlice_l113_357_3);
  assign _zz_when_ArraySlice_l113_357_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_357_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_357_4 = {1'd0, _zz_when_ArraySlice_l112_357};
  assign _zz__zz_when_ArraySlice_l173_357 = (_zz__zz_when_ArraySlice_l173_357_1 + _zz__zz_when_ArraySlice_l173_357_2);
  assign _zz__zz_when_ArraySlice_l173_357_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_357_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_357_3 = {1'd0, _zz_when_ArraySlice_l112_357};
  assign _zz_when_ArraySlice_l118_357_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_357 = _zz_when_ArraySlice_l118_357_1[5:0];
  assign _zz_when_ArraySlice_l173_357_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_357_1 = {2'd0, _zz_when_ArraySlice_l173_357_2};
  assign _zz_when_ArraySlice_l173_357_3 = (_zz_when_ArraySlice_l173_357_4 + _zz_when_ArraySlice_l173_357_8);
  assign _zz_when_ArraySlice_l173_357_4 = (_zz_when_ArraySlice_l173_357 - _zz_when_ArraySlice_l173_357_5);
  assign _zz_when_ArraySlice_l173_357_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_357_7);
  assign _zz_when_ArraySlice_l173_357_5 = {1'd0, _zz_when_ArraySlice_l173_357_6};
  assign _zz_when_ArraySlice_l173_357_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_357_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_358 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_358_1);
  assign _zz_when_ArraySlice_l165_358_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_358_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_358 = {1'd0, _zz_when_ArraySlice_l166_358_1};
  assign _zz_when_ArraySlice_l166_358_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_358_3);
  assign _zz_when_ArraySlice_l166_358_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_358_4);
  assign _zz_when_ArraySlice_l166_358_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_358 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_358 = (_zz_when_ArraySlice_l113_358_1 - _zz_when_ArraySlice_l113_358_4);
  assign _zz_when_ArraySlice_l113_358_1 = (_zz_when_ArraySlice_l113_358_2 + _zz_when_ArraySlice_l113_358_3);
  assign _zz_when_ArraySlice_l113_358_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_358_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_358_4 = {1'd0, _zz_when_ArraySlice_l112_358};
  assign _zz__zz_when_ArraySlice_l173_358 = (_zz__zz_when_ArraySlice_l173_358_1 + _zz__zz_when_ArraySlice_l173_358_2);
  assign _zz__zz_when_ArraySlice_l173_358_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_358_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_358_3 = {1'd0, _zz_when_ArraySlice_l112_358};
  assign _zz_when_ArraySlice_l118_358_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_358 = _zz_when_ArraySlice_l118_358_1[5:0];
  assign _zz_when_ArraySlice_l173_358_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_358_1 = {2'd0, _zz_when_ArraySlice_l173_358_2};
  assign _zz_when_ArraySlice_l173_358_3 = (_zz_when_ArraySlice_l173_358_4 + _zz_when_ArraySlice_l173_358_8);
  assign _zz_when_ArraySlice_l173_358_4 = (_zz_when_ArraySlice_l173_358 - _zz_when_ArraySlice_l173_358_5);
  assign _zz_when_ArraySlice_l173_358_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_358_7);
  assign _zz_when_ArraySlice_l173_358_5 = {1'd0, _zz_when_ArraySlice_l173_358_6};
  assign _zz_when_ArraySlice_l173_358_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_358_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_359 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_359_1);
  assign _zz_when_ArraySlice_l165_359_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_359_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_359 = {2'd0, _zz_when_ArraySlice_l166_359_1};
  assign _zz_when_ArraySlice_l166_359_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_359_3);
  assign _zz_when_ArraySlice_l166_359_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_359_4);
  assign _zz_when_ArraySlice_l166_359_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_359 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_359 = (_zz_when_ArraySlice_l113_359_1 - _zz_when_ArraySlice_l113_359_4);
  assign _zz_when_ArraySlice_l113_359_1 = (_zz_when_ArraySlice_l113_359_2 + _zz_when_ArraySlice_l113_359_3);
  assign _zz_when_ArraySlice_l113_359_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_359_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_359_4 = {1'd0, _zz_when_ArraySlice_l112_359};
  assign _zz__zz_when_ArraySlice_l173_359 = (_zz__zz_when_ArraySlice_l173_359_1 + _zz__zz_when_ArraySlice_l173_359_2);
  assign _zz__zz_when_ArraySlice_l173_359_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_359_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_359_3 = {1'd0, _zz_when_ArraySlice_l112_359};
  assign _zz_when_ArraySlice_l118_359_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_359 = _zz_when_ArraySlice_l118_359_1[5:0];
  assign _zz_when_ArraySlice_l173_359_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_359_1 = {3'd0, _zz_when_ArraySlice_l173_359_2};
  assign _zz_when_ArraySlice_l173_359_3 = (_zz_when_ArraySlice_l173_359_4 + _zz_when_ArraySlice_l173_359_8);
  assign _zz_when_ArraySlice_l173_359_4 = (_zz_when_ArraySlice_l173_359 - _zz_when_ArraySlice_l173_359_5);
  assign _zz_when_ArraySlice_l173_359_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_359_7);
  assign _zz_when_ArraySlice_l173_359_5 = {1'd0, _zz_when_ArraySlice_l173_359_6};
  assign _zz_when_ArraySlice_l173_359_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_359_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l268_6_1 = (_zz_when_ArraySlice_l268_6_2 + _zz_when_ArraySlice_l268_6_7);
  assign _zz_when_ArraySlice_l268_6_2 = (_zz_when_ArraySlice_l268_6_3 + _zz_when_ArraySlice_l268_6_5);
  assign _zz_when_ArraySlice_l268_6_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l268_6_4);
  assign _zz_when_ArraySlice_l268_6_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l268_6_6 = 1'b1;
  assign _zz_when_ArraySlice_l268_6_5 = {5'd0, _zz_when_ArraySlice_l268_6_6};
  assign _zz_when_ArraySlice_l268_6_7 = (bReg * 3'b110);
  assign _zz_selectReadFifo_6_47 = 1'b1;
  assign _zz_selectReadFifo_6_46 = {5'd0, _zz_selectReadFifo_6_47};
  assign _zz_when_ArraySlice_l272_6 = (_zz_when_ArraySlice_l272_6_1 % aReg);
  assign _zz_when_ArraySlice_l272_6_1 = (handshakeTimes_6_value + _zz_when_ArraySlice_l272_6_2);
  assign _zz_when_ArraySlice_l272_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l272_6_2 = {12'd0, _zz_when_ArraySlice_l272_6_3};
  assign _zz_when_ArraySlice_l276_6_1 = (selectReadFifo_6 + _zz_when_ArraySlice_l276_6_2);
  assign _zz_when_ArraySlice_l276_6_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l277_6_1 = (_zz_when_ArraySlice_l277_6_2 - _zz_when_ArraySlice_l277_6_3);
  assign _zz_when_ArraySlice_l277_6 = {7'd0, _zz_when_ArraySlice_l277_6_1};
  assign _zz_when_ArraySlice_l277_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l277_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l277_6_3 = {5'd0, _zz_when_ArraySlice_l277_6_4};
  assign _zz__zz_when_ArraySlice_l94_43 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_43 = (_zz_when_ArraySlice_l95_43_1 - _zz_when_ArraySlice_l95_43_4);
  assign _zz_when_ArraySlice_l95_43_1 = (_zz_when_ArraySlice_l95_43_2 + _zz_when_ArraySlice_l95_43_3);
  assign _zz_when_ArraySlice_l95_43_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_43_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_43_4 = {1'd0, _zz_when_ArraySlice_l94_43};
  assign _zz__zz_when_ArraySlice_l279_6 = (_zz__zz_when_ArraySlice_l279_6_1 + _zz__zz_when_ArraySlice_l279_6_2);
  assign _zz__zz_when_ArraySlice_l279_6_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l279_6_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l279_6_3 = {1'd0, _zz_when_ArraySlice_l94_43};
  assign _zz_when_ArraySlice_l99_43_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_43 = _zz_when_ArraySlice_l99_43_1[5:0];
  assign _zz_when_ArraySlice_l279_6_1 = (outSliceNumb_6_value + _zz_when_ArraySlice_l279_6_2);
  assign _zz_when_ArraySlice_l279_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l279_6_2 = {6'd0, _zz_when_ArraySlice_l279_6_3};
  assign _zz_when_ArraySlice_l279_6_4 = (_zz_when_ArraySlice_l279_6 / aReg);
  assign _zz_selectReadFifo_6_48 = (selectReadFifo_6 - _zz_selectReadFifo_6_49);
  assign _zz_selectReadFifo_6_49 = {3'd0, bReg};
  assign _zz_selectReadFifo_6_51 = 1'b1;
  assign _zz_selectReadFifo_6_50 = {5'd0, _zz_selectReadFifo_6_51};
  assign _zz_selectReadFifo_6_52 = (selectReadFifo_6 + _zz_selectReadFifo_6_53);
  assign _zz_selectReadFifo_6_53 = (3'b111 * bReg);
  assign _zz_selectReadFifo_6_55 = 1'b1;
  assign _zz_selectReadFifo_6_54 = {5'd0, _zz_selectReadFifo_6_55};
  assign _zz_when_ArraySlice_l165_360 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_360_1);
  assign _zz_when_ArraySlice_l165_360_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_360_1 = {3'd0, _zz_when_ArraySlice_l165_360_2};
  assign _zz_when_ArraySlice_l166_360 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_360_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_360_3);
  assign _zz_when_ArraySlice_l166_360_1 = {1'd0, _zz_when_ArraySlice_l166_360_2};
  assign _zz_when_ArraySlice_l166_360_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_360_4);
  assign _zz_when_ArraySlice_l166_360_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_360_4 = {3'd0, _zz_when_ArraySlice_l166_360_5};
  assign _zz__zz_when_ArraySlice_l112_360 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_360 = (_zz_when_ArraySlice_l113_360_1 - _zz_when_ArraySlice_l113_360_4);
  assign _zz_when_ArraySlice_l113_360_1 = (_zz_when_ArraySlice_l113_360_2 + _zz_when_ArraySlice_l113_360_3);
  assign _zz_when_ArraySlice_l113_360_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_360_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_360_4 = {1'd0, _zz_when_ArraySlice_l112_360};
  assign _zz__zz_when_ArraySlice_l173_360 = (_zz__zz_when_ArraySlice_l173_360_1 + _zz__zz_when_ArraySlice_l173_360_2);
  assign _zz__zz_when_ArraySlice_l173_360_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_360_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_360_3 = {1'd0, _zz_when_ArraySlice_l112_360};
  assign _zz_when_ArraySlice_l118_360_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_360 = _zz_when_ArraySlice_l118_360_1[5:0];
  assign _zz_when_ArraySlice_l173_360_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_360_2 = (_zz_when_ArraySlice_l173_360_3 + _zz_when_ArraySlice_l173_360_8);
  assign _zz_when_ArraySlice_l173_360_3 = (_zz_when_ArraySlice_l173_360 - _zz_when_ArraySlice_l173_360_4);
  assign _zz_when_ArraySlice_l173_360_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_360_6);
  assign _zz_when_ArraySlice_l173_360_4 = {1'd0, _zz_when_ArraySlice_l173_360_5};
  assign _zz_when_ArraySlice_l173_360_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_360_6 = {3'd0, _zz_when_ArraySlice_l173_360_7};
  assign _zz_when_ArraySlice_l173_360_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_361 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_361_1);
  assign _zz_when_ArraySlice_l165_361_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_361_1 = {2'd0, _zz_when_ArraySlice_l165_361_2};
  assign _zz_when_ArraySlice_l166_361 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_361_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_361_2);
  assign _zz_when_ArraySlice_l166_361_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_361_3);
  assign _zz_when_ArraySlice_l166_361_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_361_3 = {2'd0, _zz_when_ArraySlice_l166_361_4};
  assign _zz__zz_when_ArraySlice_l112_361 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_361 = (_zz_when_ArraySlice_l113_361_1 - _zz_when_ArraySlice_l113_361_4);
  assign _zz_when_ArraySlice_l113_361_1 = (_zz_when_ArraySlice_l113_361_2 + _zz_when_ArraySlice_l113_361_3);
  assign _zz_when_ArraySlice_l113_361_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_361_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_361_4 = {1'd0, _zz_when_ArraySlice_l112_361};
  assign _zz__zz_when_ArraySlice_l173_361 = (_zz__zz_when_ArraySlice_l173_361_1 + _zz__zz_when_ArraySlice_l173_361_2);
  assign _zz__zz_when_ArraySlice_l173_361_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_361_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_361_3 = {1'd0, _zz_when_ArraySlice_l112_361};
  assign _zz_when_ArraySlice_l118_361_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_361 = _zz_when_ArraySlice_l118_361_1[5:0];
  assign _zz_when_ArraySlice_l173_361_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_361_1 = {1'd0, _zz_when_ArraySlice_l173_361_2};
  assign _zz_when_ArraySlice_l173_361_3 = (_zz_when_ArraySlice_l173_361_4 + _zz_when_ArraySlice_l173_361_9);
  assign _zz_when_ArraySlice_l173_361_4 = (_zz_when_ArraySlice_l173_361 - _zz_when_ArraySlice_l173_361_5);
  assign _zz_when_ArraySlice_l173_361_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_361_7);
  assign _zz_when_ArraySlice_l173_361_5 = {1'd0, _zz_when_ArraySlice_l173_361_6};
  assign _zz_when_ArraySlice_l173_361_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_361_7 = {2'd0, _zz_when_ArraySlice_l173_361_8};
  assign _zz_when_ArraySlice_l173_361_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_362 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_362_1);
  assign _zz_when_ArraySlice_l165_362_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_362_1 = {1'd0, _zz_when_ArraySlice_l165_362_2};
  assign _zz_when_ArraySlice_l166_362 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_362_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_362_2);
  assign _zz_when_ArraySlice_l166_362_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_362_3);
  assign _zz_when_ArraySlice_l166_362_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_362_3 = {1'd0, _zz_when_ArraySlice_l166_362_4};
  assign _zz__zz_when_ArraySlice_l112_362 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_362 = (_zz_when_ArraySlice_l113_362_1 - _zz_when_ArraySlice_l113_362_4);
  assign _zz_when_ArraySlice_l113_362_1 = (_zz_when_ArraySlice_l113_362_2 + _zz_when_ArraySlice_l113_362_3);
  assign _zz_when_ArraySlice_l113_362_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_362_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_362_4 = {1'd0, _zz_when_ArraySlice_l112_362};
  assign _zz__zz_when_ArraySlice_l173_362 = (_zz__zz_when_ArraySlice_l173_362_1 + _zz__zz_when_ArraySlice_l173_362_2);
  assign _zz__zz_when_ArraySlice_l173_362_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_362_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_362_3 = {1'd0, _zz_when_ArraySlice_l112_362};
  assign _zz_when_ArraySlice_l118_362_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_362 = _zz_when_ArraySlice_l118_362_1[5:0];
  assign _zz_when_ArraySlice_l173_362_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_362_1 = {1'd0, _zz_when_ArraySlice_l173_362_2};
  assign _zz_when_ArraySlice_l173_362_3 = (_zz_when_ArraySlice_l173_362_4 + _zz_when_ArraySlice_l173_362_9);
  assign _zz_when_ArraySlice_l173_362_4 = (_zz_when_ArraySlice_l173_362 - _zz_when_ArraySlice_l173_362_5);
  assign _zz_when_ArraySlice_l173_362_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_362_7);
  assign _zz_when_ArraySlice_l173_362_5 = {1'd0, _zz_when_ArraySlice_l173_362_6};
  assign _zz_when_ArraySlice_l173_362_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_362_7 = {1'd0, _zz_when_ArraySlice_l173_362_8};
  assign _zz_when_ArraySlice_l173_362_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_363 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_363_1);
  assign _zz_when_ArraySlice_l165_363_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_363_1 = {1'd0, _zz_when_ArraySlice_l165_363_2};
  assign _zz_when_ArraySlice_l166_363 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_363_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_363_2);
  assign _zz_when_ArraySlice_l166_363_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_363_3);
  assign _zz_when_ArraySlice_l166_363_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_363_3 = {1'd0, _zz_when_ArraySlice_l166_363_4};
  assign _zz__zz_when_ArraySlice_l112_363 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_363 = (_zz_when_ArraySlice_l113_363_1 - _zz_when_ArraySlice_l113_363_4);
  assign _zz_when_ArraySlice_l113_363_1 = (_zz_when_ArraySlice_l113_363_2 + _zz_when_ArraySlice_l113_363_3);
  assign _zz_when_ArraySlice_l113_363_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_363_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_363_4 = {1'd0, _zz_when_ArraySlice_l112_363};
  assign _zz__zz_when_ArraySlice_l173_363 = (_zz__zz_when_ArraySlice_l173_363_1 + _zz__zz_when_ArraySlice_l173_363_2);
  assign _zz__zz_when_ArraySlice_l173_363_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_363_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_363_3 = {1'd0, _zz_when_ArraySlice_l112_363};
  assign _zz_when_ArraySlice_l118_363_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_363 = _zz_when_ArraySlice_l118_363_1[5:0];
  assign _zz_when_ArraySlice_l173_363_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_363_1 = {1'd0, _zz_when_ArraySlice_l173_363_2};
  assign _zz_when_ArraySlice_l173_363_3 = (_zz_when_ArraySlice_l173_363_4 + _zz_when_ArraySlice_l173_363_9);
  assign _zz_when_ArraySlice_l173_363_4 = (_zz_when_ArraySlice_l173_363 - _zz_when_ArraySlice_l173_363_5);
  assign _zz_when_ArraySlice_l173_363_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_363_7);
  assign _zz_when_ArraySlice_l173_363_5 = {1'd0, _zz_when_ArraySlice_l173_363_6};
  assign _zz_when_ArraySlice_l173_363_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_363_7 = {1'd0, _zz_when_ArraySlice_l173_363_8};
  assign _zz_when_ArraySlice_l173_363_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_364 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_364_1);
  assign _zz_when_ArraySlice_l165_364_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_364 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_364_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_364_2);
  assign _zz_when_ArraySlice_l166_364_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_364_3);
  assign _zz_when_ArraySlice_l166_364_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_364 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_364 = (_zz_when_ArraySlice_l113_364_1 - _zz_when_ArraySlice_l113_364_4);
  assign _zz_when_ArraySlice_l113_364_1 = (_zz_when_ArraySlice_l113_364_2 + _zz_when_ArraySlice_l113_364_3);
  assign _zz_when_ArraySlice_l113_364_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_364_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_364_4 = {1'd0, _zz_when_ArraySlice_l112_364};
  assign _zz__zz_when_ArraySlice_l173_364 = (_zz__zz_when_ArraySlice_l173_364_1 + _zz__zz_when_ArraySlice_l173_364_2);
  assign _zz__zz_when_ArraySlice_l173_364_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_364_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_364_3 = {1'd0, _zz_when_ArraySlice_l112_364};
  assign _zz_when_ArraySlice_l118_364_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_364 = _zz_when_ArraySlice_l118_364_1[5:0];
  assign _zz_when_ArraySlice_l173_364_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_364_1 = {1'd0, _zz_when_ArraySlice_l173_364_2};
  assign _zz_when_ArraySlice_l173_364_3 = (_zz_when_ArraySlice_l173_364_4 + _zz_when_ArraySlice_l173_364_8);
  assign _zz_when_ArraySlice_l173_364_4 = (_zz_when_ArraySlice_l173_364 - _zz_when_ArraySlice_l173_364_5);
  assign _zz_when_ArraySlice_l173_364_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_364_7);
  assign _zz_when_ArraySlice_l173_364_5 = {1'd0, _zz_when_ArraySlice_l173_364_6};
  assign _zz_when_ArraySlice_l173_364_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_364_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_365 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_365_1);
  assign _zz_when_ArraySlice_l165_365_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_365_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_365 = {1'd0, _zz_when_ArraySlice_l166_365_1};
  assign _zz_when_ArraySlice_l166_365_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_365_3);
  assign _zz_when_ArraySlice_l166_365_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_365_4);
  assign _zz_when_ArraySlice_l166_365_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_365 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_365 = (_zz_when_ArraySlice_l113_365_1 - _zz_when_ArraySlice_l113_365_4);
  assign _zz_when_ArraySlice_l113_365_1 = (_zz_when_ArraySlice_l113_365_2 + _zz_when_ArraySlice_l113_365_3);
  assign _zz_when_ArraySlice_l113_365_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_365_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_365_4 = {1'd0, _zz_when_ArraySlice_l112_365};
  assign _zz__zz_when_ArraySlice_l173_365 = (_zz__zz_when_ArraySlice_l173_365_1 + _zz__zz_when_ArraySlice_l173_365_2);
  assign _zz__zz_when_ArraySlice_l173_365_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_365_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_365_3 = {1'd0, _zz_when_ArraySlice_l112_365};
  assign _zz_when_ArraySlice_l118_365_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_365 = _zz_when_ArraySlice_l118_365_1[5:0];
  assign _zz_when_ArraySlice_l173_365_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_365_1 = {2'd0, _zz_when_ArraySlice_l173_365_2};
  assign _zz_when_ArraySlice_l173_365_3 = (_zz_when_ArraySlice_l173_365_4 + _zz_when_ArraySlice_l173_365_8);
  assign _zz_when_ArraySlice_l173_365_4 = (_zz_when_ArraySlice_l173_365 - _zz_when_ArraySlice_l173_365_5);
  assign _zz_when_ArraySlice_l173_365_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_365_7);
  assign _zz_when_ArraySlice_l173_365_5 = {1'd0, _zz_when_ArraySlice_l173_365_6};
  assign _zz_when_ArraySlice_l173_365_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_365_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_366 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_366_1);
  assign _zz_when_ArraySlice_l165_366_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_366_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_366 = {1'd0, _zz_when_ArraySlice_l166_366_1};
  assign _zz_when_ArraySlice_l166_366_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_366_3);
  assign _zz_when_ArraySlice_l166_366_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_366_4);
  assign _zz_when_ArraySlice_l166_366_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_366 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_366 = (_zz_when_ArraySlice_l113_366_1 - _zz_when_ArraySlice_l113_366_4);
  assign _zz_when_ArraySlice_l113_366_1 = (_zz_when_ArraySlice_l113_366_2 + _zz_when_ArraySlice_l113_366_3);
  assign _zz_when_ArraySlice_l113_366_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_366_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_366_4 = {1'd0, _zz_when_ArraySlice_l112_366};
  assign _zz__zz_when_ArraySlice_l173_366 = (_zz__zz_when_ArraySlice_l173_366_1 + _zz__zz_when_ArraySlice_l173_366_2);
  assign _zz__zz_when_ArraySlice_l173_366_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_366_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_366_3 = {1'd0, _zz_when_ArraySlice_l112_366};
  assign _zz_when_ArraySlice_l118_366_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_366 = _zz_when_ArraySlice_l118_366_1[5:0];
  assign _zz_when_ArraySlice_l173_366_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_366_1 = {2'd0, _zz_when_ArraySlice_l173_366_2};
  assign _zz_when_ArraySlice_l173_366_3 = (_zz_when_ArraySlice_l173_366_4 + _zz_when_ArraySlice_l173_366_8);
  assign _zz_when_ArraySlice_l173_366_4 = (_zz_when_ArraySlice_l173_366 - _zz_when_ArraySlice_l173_366_5);
  assign _zz_when_ArraySlice_l173_366_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_366_7);
  assign _zz_when_ArraySlice_l173_366_5 = {1'd0, _zz_when_ArraySlice_l173_366_6};
  assign _zz_when_ArraySlice_l173_366_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_366_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_367 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_367_1);
  assign _zz_when_ArraySlice_l165_367_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_367_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_367 = {2'd0, _zz_when_ArraySlice_l166_367_1};
  assign _zz_when_ArraySlice_l166_367_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_367_3);
  assign _zz_when_ArraySlice_l166_367_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_367_4);
  assign _zz_when_ArraySlice_l166_367_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_367 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_367 = (_zz_when_ArraySlice_l113_367_1 - _zz_when_ArraySlice_l113_367_4);
  assign _zz_when_ArraySlice_l113_367_1 = (_zz_when_ArraySlice_l113_367_2 + _zz_when_ArraySlice_l113_367_3);
  assign _zz_when_ArraySlice_l113_367_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_367_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_367_4 = {1'd0, _zz_when_ArraySlice_l112_367};
  assign _zz__zz_when_ArraySlice_l173_367 = (_zz__zz_when_ArraySlice_l173_367_1 + _zz__zz_when_ArraySlice_l173_367_2);
  assign _zz__zz_when_ArraySlice_l173_367_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_367_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_367_3 = {1'd0, _zz_when_ArraySlice_l112_367};
  assign _zz_when_ArraySlice_l118_367_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_367 = _zz_when_ArraySlice_l118_367_1[5:0];
  assign _zz_when_ArraySlice_l173_367_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_367_1 = {3'd0, _zz_when_ArraySlice_l173_367_2};
  assign _zz_when_ArraySlice_l173_367_3 = (_zz_when_ArraySlice_l173_367_4 + _zz_when_ArraySlice_l173_367_8);
  assign _zz_when_ArraySlice_l173_367_4 = (_zz_when_ArraySlice_l173_367 - _zz_when_ArraySlice_l173_367_5);
  assign _zz_when_ArraySlice_l173_367_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_367_7);
  assign _zz_when_ArraySlice_l173_367_5 = {1'd0, _zz_when_ArraySlice_l173_367_6};
  assign _zz_when_ArraySlice_l173_367_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_367_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l288_6_1 = (_zz_when_ArraySlice_l288_6_2 + _zz_when_ArraySlice_l288_6_7);
  assign _zz_when_ArraySlice_l288_6_2 = (_zz_when_ArraySlice_l288_6_3 + _zz_when_ArraySlice_l288_6_5);
  assign _zz_when_ArraySlice_l288_6_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l288_6_4);
  assign _zz_when_ArraySlice_l288_6_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_6_6 = 1'b1;
  assign _zz_when_ArraySlice_l288_6_5 = {5'd0, _zz_when_ArraySlice_l288_6_6};
  assign _zz_when_ArraySlice_l288_6_7 = (bReg * 3'b110);
  assign _zz_selectReadFifo_6_57 = 1'b1;
  assign _zz_selectReadFifo_6_56 = {5'd0, _zz_selectReadFifo_6_57};
  assign _zz_when_ArraySlice_l292_6 = (_zz_when_ArraySlice_l292_6_1 % aReg);
  assign _zz_when_ArraySlice_l292_6_1 = (handshakeTimes_6_value + _zz_when_ArraySlice_l292_6_2);
  assign _zz_when_ArraySlice_l292_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l292_6_2 = {12'd0, _zz_when_ArraySlice_l292_6_3};
  assign _zz_when_ArraySlice_l303_6_1 = (_zz_when_ArraySlice_l303_6_2 - _zz_when_ArraySlice_l303_6_3);
  assign _zz_when_ArraySlice_l303_6 = {7'd0, _zz_when_ArraySlice_l303_6_1};
  assign _zz_when_ArraySlice_l303_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l303_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l303_6_3 = {5'd0, _zz_when_ArraySlice_l303_6_4};
  assign _zz__zz_when_ArraySlice_l94_44 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_44 = (_zz_when_ArraySlice_l95_44_1 - _zz_when_ArraySlice_l95_44_4);
  assign _zz_when_ArraySlice_l95_44_1 = (_zz_when_ArraySlice_l95_44_2 + _zz_when_ArraySlice_l95_44_3);
  assign _zz_when_ArraySlice_l95_44_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_44_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_44_4 = {1'd0, _zz_when_ArraySlice_l94_44};
  assign _zz__zz_when_ArraySlice_l304_6 = (_zz__zz_when_ArraySlice_l304_6_1 + _zz__zz_when_ArraySlice_l304_6_2);
  assign _zz__zz_when_ArraySlice_l304_6_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l304_6_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l304_6_3 = {1'd0, _zz_when_ArraySlice_l94_44};
  assign _zz_when_ArraySlice_l99_44_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_44 = _zz_when_ArraySlice_l99_44_1[5:0];
  assign _zz_when_ArraySlice_l304_6_1 = (outSliceNumb_6_value + _zz_when_ArraySlice_l304_6_2);
  assign _zz_when_ArraySlice_l304_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l304_6_2 = {6'd0, _zz_when_ArraySlice_l304_6_3};
  assign _zz_when_ArraySlice_l304_6_4 = (_zz_when_ArraySlice_l304_6 / aReg);
  assign _zz_selectReadFifo_6_58 = (selectReadFifo_6 - _zz_selectReadFifo_6_59);
  assign _zz_selectReadFifo_6_59 = {3'd0, bReg};
  assign _zz_selectReadFifo_6_61 = 1'b1;
  assign _zz_selectReadFifo_6_60 = {5'd0, _zz_selectReadFifo_6_61};
  assign _zz_when_ArraySlice_l165_368 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_368_1);
  assign _zz_when_ArraySlice_l165_368_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_368_1 = {3'd0, _zz_when_ArraySlice_l165_368_2};
  assign _zz_when_ArraySlice_l166_368 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_368_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_368_3);
  assign _zz_when_ArraySlice_l166_368_1 = {1'd0, _zz_when_ArraySlice_l166_368_2};
  assign _zz_when_ArraySlice_l166_368_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_368_4);
  assign _zz_when_ArraySlice_l166_368_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_368_4 = {3'd0, _zz_when_ArraySlice_l166_368_5};
  assign _zz__zz_when_ArraySlice_l112_368 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_368 = (_zz_when_ArraySlice_l113_368_1 - _zz_when_ArraySlice_l113_368_4);
  assign _zz_when_ArraySlice_l113_368_1 = (_zz_when_ArraySlice_l113_368_2 + _zz_when_ArraySlice_l113_368_3);
  assign _zz_when_ArraySlice_l113_368_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_368_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_368_4 = {1'd0, _zz_when_ArraySlice_l112_368};
  assign _zz__zz_when_ArraySlice_l173_368 = (_zz__zz_when_ArraySlice_l173_368_1 + _zz__zz_when_ArraySlice_l173_368_2);
  assign _zz__zz_when_ArraySlice_l173_368_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_368_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_368_3 = {1'd0, _zz_when_ArraySlice_l112_368};
  assign _zz_when_ArraySlice_l118_368_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_368 = _zz_when_ArraySlice_l118_368_1[5:0];
  assign _zz_when_ArraySlice_l173_368_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_368_2 = (_zz_when_ArraySlice_l173_368_3 + _zz_when_ArraySlice_l173_368_8);
  assign _zz_when_ArraySlice_l173_368_3 = (_zz_when_ArraySlice_l173_368 - _zz_when_ArraySlice_l173_368_4);
  assign _zz_when_ArraySlice_l173_368_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_368_6);
  assign _zz_when_ArraySlice_l173_368_4 = {1'd0, _zz_when_ArraySlice_l173_368_5};
  assign _zz_when_ArraySlice_l173_368_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_368_6 = {3'd0, _zz_when_ArraySlice_l173_368_7};
  assign _zz_when_ArraySlice_l173_368_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_369 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_369_1);
  assign _zz_when_ArraySlice_l165_369_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_369_1 = {2'd0, _zz_when_ArraySlice_l165_369_2};
  assign _zz_when_ArraySlice_l166_369 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_369_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_369_2);
  assign _zz_when_ArraySlice_l166_369_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_369_3);
  assign _zz_when_ArraySlice_l166_369_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_369_3 = {2'd0, _zz_when_ArraySlice_l166_369_4};
  assign _zz__zz_when_ArraySlice_l112_369 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_369 = (_zz_when_ArraySlice_l113_369_1 - _zz_when_ArraySlice_l113_369_4);
  assign _zz_when_ArraySlice_l113_369_1 = (_zz_when_ArraySlice_l113_369_2 + _zz_when_ArraySlice_l113_369_3);
  assign _zz_when_ArraySlice_l113_369_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_369_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_369_4 = {1'd0, _zz_when_ArraySlice_l112_369};
  assign _zz__zz_when_ArraySlice_l173_369 = (_zz__zz_when_ArraySlice_l173_369_1 + _zz__zz_when_ArraySlice_l173_369_2);
  assign _zz__zz_when_ArraySlice_l173_369_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_369_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_369_3 = {1'd0, _zz_when_ArraySlice_l112_369};
  assign _zz_when_ArraySlice_l118_369_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_369 = _zz_when_ArraySlice_l118_369_1[5:0];
  assign _zz_when_ArraySlice_l173_369_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_369_1 = {1'd0, _zz_when_ArraySlice_l173_369_2};
  assign _zz_when_ArraySlice_l173_369_3 = (_zz_when_ArraySlice_l173_369_4 + _zz_when_ArraySlice_l173_369_9);
  assign _zz_when_ArraySlice_l173_369_4 = (_zz_when_ArraySlice_l173_369 - _zz_when_ArraySlice_l173_369_5);
  assign _zz_when_ArraySlice_l173_369_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_369_7);
  assign _zz_when_ArraySlice_l173_369_5 = {1'd0, _zz_when_ArraySlice_l173_369_6};
  assign _zz_when_ArraySlice_l173_369_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_369_7 = {2'd0, _zz_when_ArraySlice_l173_369_8};
  assign _zz_when_ArraySlice_l173_369_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_370 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_370_1);
  assign _zz_when_ArraySlice_l165_370_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_370_1 = {1'd0, _zz_when_ArraySlice_l165_370_2};
  assign _zz_when_ArraySlice_l166_370 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_370_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_370_2);
  assign _zz_when_ArraySlice_l166_370_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_370_3);
  assign _zz_when_ArraySlice_l166_370_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_370_3 = {1'd0, _zz_when_ArraySlice_l166_370_4};
  assign _zz__zz_when_ArraySlice_l112_370 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_370 = (_zz_when_ArraySlice_l113_370_1 - _zz_when_ArraySlice_l113_370_4);
  assign _zz_when_ArraySlice_l113_370_1 = (_zz_when_ArraySlice_l113_370_2 + _zz_when_ArraySlice_l113_370_3);
  assign _zz_when_ArraySlice_l113_370_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_370_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_370_4 = {1'd0, _zz_when_ArraySlice_l112_370};
  assign _zz__zz_when_ArraySlice_l173_370 = (_zz__zz_when_ArraySlice_l173_370_1 + _zz__zz_when_ArraySlice_l173_370_2);
  assign _zz__zz_when_ArraySlice_l173_370_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_370_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_370_3 = {1'd0, _zz_when_ArraySlice_l112_370};
  assign _zz_when_ArraySlice_l118_370_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_370 = _zz_when_ArraySlice_l118_370_1[5:0];
  assign _zz_when_ArraySlice_l173_370_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_370_1 = {1'd0, _zz_when_ArraySlice_l173_370_2};
  assign _zz_when_ArraySlice_l173_370_3 = (_zz_when_ArraySlice_l173_370_4 + _zz_when_ArraySlice_l173_370_9);
  assign _zz_when_ArraySlice_l173_370_4 = (_zz_when_ArraySlice_l173_370 - _zz_when_ArraySlice_l173_370_5);
  assign _zz_when_ArraySlice_l173_370_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_370_7);
  assign _zz_when_ArraySlice_l173_370_5 = {1'd0, _zz_when_ArraySlice_l173_370_6};
  assign _zz_when_ArraySlice_l173_370_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_370_7 = {1'd0, _zz_when_ArraySlice_l173_370_8};
  assign _zz_when_ArraySlice_l173_370_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_371 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_371_1);
  assign _zz_when_ArraySlice_l165_371_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_371_1 = {1'd0, _zz_when_ArraySlice_l165_371_2};
  assign _zz_when_ArraySlice_l166_371 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_371_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_371_2);
  assign _zz_when_ArraySlice_l166_371_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_371_3);
  assign _zz_when_ArraySlice_l166_371_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_371_3 = {1'd0, _zz_when_ArraySlice_l166_371_4};
  assign _zz__zz_when_ArraySlice_l112_371 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_371 = (_zz_when_ArraySlice_l113_371_1 - _zz_when_ArraySlice_l113_371_4);
  assign _zz_when_ArraySlice_l113_371_1 = (_zz_when_ArraySlice_l113_371_2 + _zz_when_ArraySlice_l113_371_3);
  assign _zz_when_ArraySlice_l113_371_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_371_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_371_4 = {1'd0, _zz_when_ArraySlice_l112_371};
  assign _zz__zz_when_ArraySlice_l173_371 = (_zz__zz_when_ArraySlice_l173_371_1 + _zz__zz_when_ArraySlice_l173_371_2);
  assign _zz__zz_when_ArraySlice_l173_371_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_371_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_371_3 = {1'd0, _zz_when_ArraySlice_l112_371};
  assign _zz_when_ArraySlice_l118_371_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_371 = _zz_when_ArraySlice_l118_371_1[5:0];
  assign _zz_when_ArraySlice_l173_371_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_371_1 = {1'd0, _zz_when_ArraySlice_l173_371_2};
  assign _zz_when_ArraySlice_l173_371_3 = (_zz_when_ArraySlice_l173_371_4 + _zz_when_ArraySlice_l173_371_9);
  assign _zz_when_ArraySlice_l173_371_4 = (_zz_when_ArraySlice_l173_371 - _zz_when_ArraySlice_l173_371_5);
  assign _zz_when_ArraySlice_l173_371_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_371_7);
  assign _zz_when_ArraySlice_l173_371_5 = {1'd0, _zz_when_ArraySlice_l173_371_6};
  assign _zz_when_ArraySlice_l173_371_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_371_7 = {1'd0, _zz_when_ArraySlice_l173_371_8};
  assign _zz_when_ArraySlice_l173_371_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_372 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_372_1);
  assign _zz_when_ArraySlice_l165_372_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_372 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_372_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_372_2);
  assign _zz_when_ArraySlice_l166_372_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_372_3);
  assign _zz_when_ArraySlice_l166_372_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_372 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_372 = (_zz_when_ArraySlice_l113_372_1 - _zz_when_ArraySlice_l113_372_4);
  assign _zz_when_ArraySlice_l113_372_1 = (_zz_when_ArraySlice_l113_372_2 + _zz_when_ArraySlice_l113_372_3);
  assign _zz_when_ArraySlice_l113_372_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_372_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_372_4 = {1'd0, _zz_when_ArraySlice_l112_372};
  assign _zz__zz_when_ArraySlice_l173_372 = (_zz__zz_when_ArraySlice_l173_372_1 + _zz__zz_when_ArraySlice_l173_372_2);
  assign _zz__zz_when_ArraySlice_l173_372_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_372_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_372_3 = {1'd0, _zz_when_ArraySlice_l112_372};
  assign _zz_when_ArraySlice_l118_372_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_372 = _zz_when_ArraySlice_l118_372_1[5:0];
  assign _zz_when_ArraySlice_l173_372_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_372_1 = {1'd0, _zz_when_ArraySlice_l173_372_2};
  assign _zz_when_ArraySlice_l173_372_3 = (_zz_when_ArraySlice_l173_372_4 + _zz_when_ArraySlice_l173_372_8);
  assign _zz_when_ArraySlice_l173_372_4 = (_zz_when_ArraySlice_l173_372 - _zz_when_ArraySlice_l173_372_5);
  assign _zz_when_ArraySlice_l173_372_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_372_7);
  assign _zz_when_ArraySlice_l173_372_5 = {1'd0, _zz_when_ArraySlice_l173_372_6};
  assign _zz_when_ArraySlice_l173_372_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_372_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_373 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_373_1);
  assign _zz_when_ArraySlice_l165_373_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_373_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_373 = {1'd0, _zz_when_ArraySlice_l166_373_1};
  assign _zz_when_ArraySlice_l166_373_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_373_3);
  assign _zz_when_ArraySlice_l166_373_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_373_4);
  assign _zz_when_ArraySlice_l166_373_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_373 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_373 = (_zz_when_ArraySlice_l113_373_1 - _zz_when_ArraySlice_l113_373_4);
  assign _zz_when_ArraySlice_l113_373_1 = (_zz_when_ArraySlice_l113_373_2 + _zz_when_ArraySlice_l113_373_3);
  assign _zz_when_ArraySlice_l113_373_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_373_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_373_4 = {1'd0, _zz_when_ArraySlice_l112_373};
  assign _zz__zz_when_ArraySlice_l173_373 = (_zz__zz_when_ArraySlice_l173_373_1 + _zz__zz_when_ArraySlice_l173_373_2);
  assign _zz__zz_when_ArraySlice_l173_373_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_373_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_373_3 = {1'd0, _zz_when_ArraySlice_l112_373};
  assign _zz_when_ArraySlice_l118_373_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_373 = _zz_when_ArraySlice_l118_373_1[5:0];
  assign _zz_when_ArraySlice_l173_373_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_373_1 = {2'd0, _zz_when_ArraySlice_l173_373_2};
  assign _zz_when_ArraySlice_l173_373_3 = (_zz_when_ArraySlice_l173_373_4 + _zz_when_ArraySlice_l173_373_8);
  assign _zz_when_ArraySlice_l173_373_4 = (_zz_when_ArraySlice_l173_373 - _zz_when_ArraySlice_l173_373_5);
  assign _zz_when_ArraySlice_l173_373_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_373_7);
  assign _zz_when_ArraySlice_l173_373_5 = {1'd0, _zz_when_ArraySlice_l173_373_6};
  assign _zz_when_ArraySlice_l173_373_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_373_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_374 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_374_1);
  assign _zz_when_ArraySlice_l165_374_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_374_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_374 = {1'd0, _zz_when_ArraySlice_l166_374_1};
  assign _zz_when_ArraySlice_l166_374_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_374_3);
  assign _zz_when_ArraySlice_l166_374_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_374_4);
  assign _zz_when_ArraySlice_l166_374_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_374 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_374 = (_zz_when_ArraySlice_l113_374_1 - _zz_when_ArraySlice_l113_374_4);
  assign _zz_when_ArraySlice_l113_374_1 = (_zz_when_ArraySlice_l113_374_2 + _zz_when_ArraySlice_l113_374_3);
  assign _zz_when_ArraySlice_l113_374_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_374_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_374_4 = {1'd0, _zz_when_ArraySlice_l112_374};
  assign _zz__zz_when_ArraySlice_l173_374 = (_zz__zz_when_ArraySlice_l173_374_1 + _zz__zz_when_ArraySlice_l173_374_2);
  assign _zz__zz_when_ArraySlice_l173_374_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_374_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_374_3 = {1'd0, _zz_when_ArraySlice_l112_374};
  assign _zz_when_ArraySlice_l118_374_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_374 = _zz_when_ArraySlice_l118_374_1[5:0];
  assign _zz_when_ArraySlice_l173_374_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_374_1 = {2'd0, _zz_when_ArraySlice_l173_374_2};
  assign _zz_when_ArraySlice_l173_374_3 = (_zz_when_ArraySlice_l173_374_4 + _zz_when_ArraySlice_l173_374_8);
  assign _zz_when_ArraySlice_l173_374_4 = (_zz_when_ArraySlice_l173_374 - _zz_when_ArraySlice_l173_374_5);
  assign _zz_when_ArraySlice_l173_374_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_374_7);
  assign _zz_when_ArraySlice_l173_374_5 = {1'd0, _zz_when_ArraySlice_l173_374_6};
  assign _zz_when_ArraySlice_l173_374_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_374_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_375 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_375_1);
  assign _zz_when_ArraySlice_l165_375_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_375_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_375 = {2'd0, _zz_when_ArraySlice_l166_375_1};
  assign _zz_when_ArraySlice_l166_375_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_375_3);
  assign _zz_when_ArraySlice_l166_375_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_375_4);
  assign _zz_when_ArraySlice_l166_375_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_375 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_375 = (_zz_when_ArraySlice_l113_375_1 - _zz_when_ArraySlice_l113_375_4);
  assign _zz_when_ArraySlice_l113_375_1 = (_zz_when_ArraySlice_l113_375_2 + _zz_when_ArraySlice_l113_375_3);
  assign _zz_when_ArraySlice_l113_375_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_375_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_375_4 = {1'd0, _zz_when_ArraySlice_l112_375};
  assign _zz__zz_when_ArraySlice_l173_375 = (_zz__zz_when_ArraySlice_l173_375_1 + _zz__zz_when_ArraySlice_l173_375_2);
  assign _zz__zz_when_ArraySlice_l173_375_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_375_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_375_3 = {1'd0, _zz_when_ArraySlice_l112_375};
  assign _zz_when_ArraySlice_l118_375_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_375 = _zz_when_ArraySlice_l118_375_1[5:0];
  assign _zz_when_ArraySlice_l173_375_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_375_1 = {3'd0, _zz_when_ArraySlice_l173_375_2};
  assign _zz_when_ArraySlice_l173_375_3 = (_zz_when_ArraySlice_l173_375_4 + _zz_when_ArraySlice_l173_375_8);
  assign _zz_when_ArraySlice_l173_375_4 = (_zz_when_ArraySlice_l173_375 - _zz_when_ArraySlice_l173_375_5);
  assign _zz_when_ArraySlice_l173_375_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_375_7);
  assign _zz_when_ArraySlice_l173_375_5 = {1'd0, _zz_when_ArraySlice_l173_375_6};
  assign _zz_when_ArraySlice_l173_375_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_375_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_6_63 = 1'b1;
  assign _zz_selectReadFifo_6_62 = {5'd0, _zz_selectReadFifo_6_63};
  assign _zz_when_ArraySlice_l315_6 = (_zz_when_ArraySlice_l315_6_1 % aReg);
  assign _zz_when_ArraySlice_l315_6_1 = (handshakeTimes_6_value + _zz_when_ArraySlice_l315_6_2);
  assign _zz_when_ArraySlice_l315_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l315_6_2 = {12'd0, _zz_when_ArraySlice_l315_6_3};
  assign _zz_when_ArraySlice_l301_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l301_6_1);
  assign _zz_when_ArraySlice_l301_6_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l322_6_1 = (_zz_when_ArraySlice_l322_6_2 - _zz_when_ArraySlice_l322_6_3);
  assign _zz_when_ArraySlice_l322_6 = {7'd0, _zz_when_ArraySlice_l322_6_1};
  assign _zz_when_ArraySlice_l322_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l322_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l322_6_3 = {5'd0, _zz_when_ArraySlice_l322_6_4};
  assign _zz_when_ArraySlice_l240_7 = (selectReadFifo_7 + _zz_when_ArraySlice_l240_7_1);
  assign _zz_when_ArraySlice_l240_7_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l241_7_1 = (selectReadFifo_7 + _zz_when_ArraySlice_l241_7_2);
  assign _zz_when_ArraySlice_l241_7_2 = (bReg * 3'b111);
  assign _zz__zz_outputStreamArrayData_7_valid_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l247_7_1 = 1'b1;
  assign _zz_when_ArraySlice_l247_7 = {6'd0, _zz_when_ArraySlice_l247_7_1};
  assign _zz_when_ArraySlice_l247_7_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l247_7_4);
  assign _zz_when_ArraySlice_l247_7_4 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l248_7_1 = (_zz_when_ArraySlice_l248_7_2 - _zz_when_ArraySlice_l248_7_3);
  assign _zz_when_ArraySlice_l248_7 = {7'd0, _zz_when_ArraySlice_l248_7_1};
  assign _zz_when_ArraySlice_l248_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l248_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l248_7_3 = {5'd0, _zz_when_ArraySlice_l248_7_4};
  assign _zz_selectReadFifo_7_32 = (selectReadFifo_7 - _zz_selectReadFifo_7_33);
  assign _zz_selectReadFifo_7_33 = {3'd0, bReg};
  assign _zz_selectReadFifo_7_35 = 1'b1;
  assign _zz_selectReadFifo_7_34 = {5'd0, _zz_selectReadFifo_7_35};
  assign _zz_selectReadFifo_7_37 = 1'b1;
  assign _zz_selectReadFifo_7_36 = {5'd0, _zz_selectReadFifo_7_37};
  assign _zz_when_ArraySlice_l251_7 = (_zz_when_ArraySlice_l251_7_1 % aReg);
  assign _zz_when_ArraySlice_l251_7_1 = (handshakeTimes_7_value + _zz_when_ArraySlice_l251_7_2);
  assign _zz_when_ArraySlice_l251_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l251_7_2 = {12'd0, _zz_when_ArraySlice_l251_7_3};
  assign _zz_when_ArraySlice_l256_7_1 = (selectReadFifo_7 + _zz_when_ArraySlice_l256_7_2);
  assign _zz_when_ArraySlice_l256_7_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l256_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l256_7_3 = {6'd0, _zz_when_ArraySlice_l256_7_4};
  assign _zz_when_ArraySlice_l257_7_1 = (_zz_when_ArraySlice_l257_7_2 - _zz_when_ArraySlice_l257_7_3);
  assign _zz_when_ArraySlice_l257_7 = {7'd0, _zz_when_ArraySlice_l257_7_1};
  assign _zz_when_ArraySlice_l257_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l257_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l257_7_3 = {5'd0, _zz_when_ArraySlice_l257_7_4};
  assign _zz__zz_when_ArraySlice_l94_45 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_45 = (_zz_when_ArraySlice_l95_45_1 - _zz_when_ArraySlice_l95_45_4);
  assign _zz_when_ArraySlice_l95_45_1 = (_zz_when_ArraySlice_l95_45_2 + _zz_when_ArraySlice_l95_45_3);
  assign _zz_when_ArraySlice_l95_45_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_45_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_45_4 = {1'd0, _zz_when_ArraySlice_l94_45};
  assign _zz__zz_when_ArraySlice_l259_7 = (_zz__zz_when_ArraySlice_l259_7_1 + _zz__zz_when_ArraySlice_l259_7_2);
  assign _zz__zz_when_ArraySlice_l259_7_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l259_7_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l259_7_3 = {1'd0, _zz_when_ArraySlice_l94_45};
  assign _zz_when_ArraySlice_l99_45_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_45 = _zz_when_ArraySlice_l99_45_1[5:0];
  assign _zz_when_ArraySlice_l259_7_1 = (outSliceNumb_7_value + _zz_when_ArraySlice_l259_7_2);
  assign _zz_when_ArraySlice_l259_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l259_7_2 = {6'd0, _zz_when_ArraySlice_l259_7_3};
  assign _zz_when_ArraySlice_l259_7_4 = (_zz_when_ArraySlice_l259_7 / aReg);
  assign _zz_selectReadFifo_7_38 = (selectReadFifo_7 - _zz_selectReadFifo_7_39);
  assign _zz_selectReadFifo_7_39 = {3'd0, bReg};
  assign _zz_selectReadFifo_7_41 = 1'b1;
  assign _zz_selectReadFifo_7_40 = {5'd0, _zz_selectReadFifo_7_41};
  assign _zz_selectReadFifo_7_42 = (selectReadFifo_7 + _zz_selectReadFifo_7_43);
  assign _zz_selectReadFifo_7_43 = (3'b111 * bReg);
  assign _zz_selectReadFifo_7_45 = 1'b1;
  assign _zz_selectReadFifo_7_44 = {5'd0, _zz_selectReadFifo_7_45};
  assign _zz_when_ArraySlice_l165_376 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_376_1);
  assign _zz_when_ArraySlice_l165_376_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_376_1 = {3'd0, _zz_when_ArraySlice_l165_376_2};
  assign _zz_when_ArraySlice_l166_376 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_376_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_376_3);
  assign _zz_when_ArraySlice_l166_376_1 = {1'd0, _zz_when_ArraySlice_l166_376_2};
  assign _zz_when_ArraySlice_l166_376_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_376_4);
  assign _zz_when_ArraySlice_l166_376_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_376_4 = {3'd0, _zz_when_ArraySlice_l166_376_5};
  assign _zz__zz_when_ArraySlice_l112_376 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_376 = (_zz_when_ArraySlice_l113_376_1 - _zz_when_ArraySlice_l113_376_4);
  assign _zz_when_ArraySlice_l113_376_1 = (_zz_when_ArraySlice_l113_376_2 + _zz_when_ArraySlice_l113_376_3);
  assign _zz_when_ArraySlice_l113_376_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_376_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_376_4 = {1'd0, _zz_when_ArraySlice_l112_376};
  assign _zz__zz_when_ArraySlice_l173_376 = (_zz__zz_when_ArraySlice_l173_376_1 + _zz__zz_when_ArraySlice_l173_376_2);
  assign _zz__zz_when_ArraySlice_l173_376_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_376_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_376_3 = {1'd0, _zz_when_ArraySlice_l112_376};
  assign _zz_when_ArraySlice_l118_376_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_376 = _zz_when_ArraySlice_l118_376_1[5:0];
  assign _zz_when_ArraySlice_l173_376_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_376_2 = (_zz_when_ArraySlice_l173_376_3 + _zz_when_ArraySlice_l173_376_8);
  assign _zz_when_ArraySlice_l173_376_3 = (_zz_when_ArraySlice_l173_376 - _zz_when_ArraySlice_l173_376_4);
  assign _zz_when_ArraySlice_l173_376_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_376_6);
  assign _zz_when_ArraySlice_l173_376_4 = {1'd0, _zz_when_ArraySlice_l173_376_5};
  assign _zz_when_ArraySlice_l173_376_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_376_6 = {3'd0, _zz_when_ArraySlice_l173_376_7};
  assign _zz_when_ArraySlice_l173_376_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_377 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_377_1);
  assign _zz_when_ArraySlice_l165_377_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_377_1 = {2'd0, _zz_when_ArraySlice_l165_377_2};
  assign _zz_when_ArraySlice_l166_377 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_377_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_377_2);
  assign _zz_when_ArraySlice_l166_377_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_377_3);
  assign _zz_when_ArraySlice_l166_377_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_377_3 = {2'd0, _zz_when_ArraySlice_l166_377_4};
  assign _zz__zz_when_ArraySlice_l112_377 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_377 = (_zz_when_ArraySlice_l113_377_1 - _zz_when_ArraySlice_l113_377_4);
  assign _zz_when_ArraySlice_l113_377_1 = (_zz_when_ArraySlice_l113_377_2 + _zz_when_ArraySlice_l113_377_3);
  assign _zz_when_ArraySlice_l113_377_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_377_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_377_4 = {1'd0, _zz_when_ArraySlice_l112_377};
  assign _zz__zz_when_ArraySlice_l173_377 = (_zz__zz_when_ArraySlice_l173_377_1 + _zz__zz_when_ArraySlice_l173_377_2);
  assign _zz__zz_when_ArraySlice_l173_377_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_377_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_377_3 = {1'd0, _zz_when_ArraySlice_l112_377};
  assign _zz_when_ArraySlice_l118_377_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_377 = _zz_when_ArraySlice_l118_377_1[5:0];
  assign _zz_when_ArraySlice_l173_377_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_377_1 = {1'd0, _zz_when_ArraySlice_l173_377_2};
  assign _zz_when_ArraySlice_l173_377_3 = (_zz_when_ArraySlice_l173_377_4 + _zz_when_ArraySlice_l173_377_9);
  assign _zz_when_ArraySlice_l173_377_4 = (_zz_when_ArraySlice_l173_377 - _zz_when_ArraySlice_l173_377_5);
  assign _zz_when_ArraySlice_l173_377_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_377_7);
  assign _zz_when_ArraySlice_l173_377_5 = {1'd0, _zz_when_ArraySlice_l173_377_6};
  assign _zz_when_ArraySlice_l173_377_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_377_7 = {2'd0, _zz_when_ArraySlice_l173_377_8};
  assign _zz_when_ArraySlice_l173_377_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_378 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_378_1);
  assign _zz_when_ArraySlice_l165_378_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_378_1 = {1'd0, _zz_when_ArraySlice_l165_378_2};
  assign _zz_when_ArraySlice_l166_378 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_378_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_378_2);
  assign _zz_when_ArraySlice_l166_378_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_378_3);
  assign _zz_when_ArraySlice_l166_378_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_378_3 = {1'd0, _zz_when_ArraySlice_l166_378_4};
  assign _zz__zz_when_ArraySlice_l112_378 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_378 = (_zz_when_ArraySlice_l113_378_1 - _zz_when_ArraySlice_l113_378_4);
  assign _zz_when_ArraySlice_l113_378_1 = (_zz_when_ArraySlice_l113_378_2 + _zz_when_ArraySlice_l113_378_3);
  assign _zz_when_ArraySlice_l113_378_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_378_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_378_4 = {1'd0, _zz_when_ArraySlice_l112_378};
  assign _zz__zz_when_ArraySlice_l173_378 = (_zz__zz_when_ArraySlice_l173_378_1 + _zz__zz_when_ArraySlice_l173_378_2);
  assign _zz__zz_when_ArraySlice_l173_378_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_378_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_378_3 = {1'd0, _zz_when_ArraySlice_l112_378};
  assign _zz_when_ArraySlice_l118_378_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_378 = _zz_when_ArraySlice_l118_378_1[5:0];
  assign _zz_when_ArraySlice_l173_378_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_378_1 = {1'd0, _zz_when_ArraySlice_l173_378_2};
  assign _zz_when_ArraySlice_l173_378_3 = (_zz_when_ArraySlice_l173_378_4 + _zz_when_ArraySlice_l173_378_9);
  assign _zz_when_ArraySlice_l173_378_4 = (_zz_when_ArraySlice_l173_378 - _zz_when_ArraySlice_l173_378_5);
  assign _zz_when_ArraySlice_l173_378_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_378_7);
  assign _zz_when_ArraySlice_l173_378_5 = {1'd0, _zz_when_ArraySlice_l173_378_6};
  assign _zz_when_ArraySlice_l173_378_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_378_7 = {1'd0, _zz_when_ArraySlice_l173_378_8};
  assign _zz_when_ArraySlice_l173_378_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_379 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_379_1);
  assign _zz_when_ArraySlice_l165_379_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_379_1 = {1'd0, _zz_when_ArraySlice_l165_379_2};
  assign _zz_when_ArraySlice_l166_379 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_379_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_379_2);
  assign _zz_when_ArraySlice_l166_379_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_379_3);
  assign _zz_when_ArraySlice_l166_379_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_379_3 = {1'd0, _zz_when_ArraySlice_l166_379_4};
  assign _zz__zz_when_ArraySlice_l112_379 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_379 = (_zz_when_ArraySlice_l113_379_1 - _zz_when_ArraySlice_l113_379_4);
  assign _zz_when_ArraySlice_l113_379_1 = (_zz_when_ArraySlice_l113_379_2 + _zz_when_ArraySlice_l113_379_3);
  assign _zz_when_ArraySlice_l113_379_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_379_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_379_4 = {1'd0, _zz_when_ArraySlice_l112_379};
  assign _zz__zz_when_ArraySlice_l173_379 = (_zz__zz_when_ArraySlice_l173_379_1 + _zz__zz_when_ArraySlice_l173_379_2);
  assign _zz__zz_when_ArraySlice_l173_379_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_379_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_379_3 = {1'd0, _zz_when_ArraySlice_l112_379};
  assign _zz_when_ArraySlice_l118_379_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_379 = _zz_when_ArraySlice_l118_379_1[5:0];
  assign _zz_when_ArraySlice_l173_379_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_379_1 = {1'd0, _zz_when_ArraySlice_l173_379_2};
  assign _zz_when_ArraySlice_l173_379_3 = (_zz_when_ArraySlice_l173_379_4 + _zz_when_ArraySlice_l173_379_9);
  assign _zz_when_ArraySlice_l173_379_4 = (_zz_when_ArraySlice_l173_379 - _zz_when_ArraySlice_l173_379_5);
  assign _zz_when_ArraySlice_l173_379_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_379_7);
  assign _zz_when_ArraySlice_l173_379_5 = {1'd0, _zz_when_ArraySlice_l173_379_6};
  assign _zz_when_ArraySlice_l173_379_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_379_7 = {1'd0, _zz_when_ArraySlice_l173_379_8};
  assign _zz_when_ArraySlice_l173_379_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_380 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_380_1);
  assign _zz_when_ArraySlice_l165_380_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_380 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_380_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_380_2);
  assign _zz_when_ArraySlice_l166_380_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_380_3);
  assign _zz_when_ArraySlice_l166_380_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_380 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_380 = (_zz_when_ArraySlice_l113_380_1 - _zz_when_ArraySlice_l113_380_4);
  assign _zz_when_ArraySlice_l113_380_1 = (_zz_when_ArraySlice_l113_380_2 + _zz_when_ArraySlice_l113_380_3);
  assign _zz_when_ArraySlice_l113_380_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_380_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_380_4 = {1'd0, _zz_when_ArraySlice_l112_380};
  assign _zz__zz_when_ArraySlice_l173_380 = (_zz__zz_when_ArraySlice_l173_380_1 + _zz__zz_when_ArraySlice_l173_380_2);
  assign _zz__zz_when_ArraySlice_l173_380_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_380_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_380_3 = {1'd0, _zz_when_ArraySlice_l112_380};
  assign _zz_when_ArraySlice_l118_380_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_380 = _zz_when_ArraySlice_l118_380_1[5:0];
  assign _zz_when_ArraySlice_l173_380_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_380_1 = {1'd0, _zz_when_ArraySlice_l173_380_2};
  assign _zz_when_ArraySlice_l173_380_3 = (_zz_when_ArraySlice_l173_380_4 + _zz_when_ArraySlice_l173_380_8);
  assign _zz_when_ArraySlice_l173_380_4 = (_zz_when_ArraySlice_l173_380 - _zz_when_ArraySlice_l173_380_5);
  assign _zz_when_ArraySlice_l173_380_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_380_7);
  assign _zz_when_ArraySlice_l173_380_5 = {1'd0, _zz_when_ArraySlice_l173_380_6};
  assign _zz_when_ArraySlice_l173_380_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_380_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_381 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_381_1);
  assign _zz_when_ArraySlice_l165_381_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_381_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_381 = {1'd0, _zz_when_ArraySlice_l166_381_1};
  assign _zz_when_ArraySlice_l166_381_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_381_3);
  assign _zz_when_ArraySlice_l166_381_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_381_4);
  assign _zz_when_ArraySlice_l166_381_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_381 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_381 = (_zz_when_ArraySlice_l113_381_1 - _zz_when_ArraySlice_l113_381_4);
  assign _zz_when_ArraySlice_l113_381_1 = (_zz_when_ArraySlice_l113_381_2 + _zz_when_ArraySlice_l113_381_3);
  assign _zz_when_ArraySlice_l113_381_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_381_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_381_4 = {1'd0, _zz_when_ArraySlice_l112_381};
  assign _zz__zz_when_ArraySlice_l173_381 = (_zz__zz_when_ArraySlice_l173_381_1 + _zz__zz_when_ArraySlice_l173_381_2);
  assign _zz__zz_when_ArraySlice_l173_381_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_381_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_381_3 = {1'd0, _zz_when_ArraySlice_l112_381};
  assign _zz_when_ArraySlice_l118_381_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_381 = _zz_when_ArraySlice_l118_381_1[5:0];
  assign _zz_when_ArraySlice_l173_381_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_381_1 = {2'd0, _zz_when_ArraySlice_l173_381_2};
  assign _zz_when_ArraySlice_l173_381_3 = (_zz_when_ArraySlice_l173_381_4 + _zz_when_ArraySlice_l173_381_8);
  assign _zz_when_ArraySlice_l173_381_4 = (_zz_when_ArraySlice_l173_381 - _zz_when_ArraySlice_l173_381_5);
  assign _zz_when_ArraySlice_l173_381_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_381_7);
  assign _zz_when_ArraySlice_l173_381_5 = {1'd0, _zz_when_ArraySlice_l173_381_6};
  assign _zz_when_ArraySlice_l173_381_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_381_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_382 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_382_1);
  assign _zz_when_ArraySlice_l165_382_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_382_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_382 = {1'd0, _zz_when_ArraySlice_l166_382_1};
  assign _zz_when_ArraySlice_l166_382_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_382_3);
  assign _zz_when_ArraySlice_l166_382_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_382_4);
  assign _zz_when_ArraySlice_l166_382_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_382 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_382 = (_zz_when_ArraySlice_l113_382_1 - _zz_when_ArraySlice_l113_382_4);
  assign _zz_when_ArraySlice_l113_382_1 = (_zz_when_ArraySlice_l113_382_2 + _zz_when_ArraySlice_l113_382_3);
  assign _zz_when_ArraySlice_l113_382_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_382_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_382_4 = {1'd0, _zz_when_ArraySlice_l112_382};
  assign _zz__zz_when_ArraySlice_l173_382 = (_zz__zz_when_ArraySlice_l173_382_1 + _zz__zz_when_ArraySlice_l173_382_2);
  assign _zz__zz_when_ArraySlice_l173_382_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_382_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_382_3 = {1'd0, _zz_when_ArraySlice_l112_382};
  assign _zz_when_ArraySlice_l118_382_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_382 = _zz_when_ArraySlice_l118_382_1[5:0];
  assign _zz_when_ArraySlice_l173_382_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_382_1 = {2'd0, _zz_when_ArraySlice_l173_382_2};
  assign _zz_when_ArraySlice_l173_382_3 = (_zz_when_ArraySlice_l173_382_4 + _zz_when_ArraySlice_l173_382_8);
  assign _zz_when_ArraySlice_l173_382_4 = (_zz_when_ArraySlice_l173_382 - _zz_when_ArraySlice_l173_382_5);
  assign _zz_when_ArraySlice_l173_382_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_382_7);
  assign _zz_when_ArraySlice_l173_382_5 = {1'd0, _zz_when_ArraySlice_l173_382_6};
  assign _zz_when_ArraySlice_l173_382_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_382_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_383 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_383_1);
  assign _zz_when_ArraySlice_l165_383_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_383_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_383 = {2'd0, _zz_when_ArraySlice_l166_383_1};
  assign _zz_when_ArraySlice_l166_383_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_383_3);
  assign _zz_when_ArraySlice_l166_383_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_383_4);
  assign _zz_when_ArraySlice_l166_383_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_383 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_383 = (_zz_when_ArraySlice_l113_383_1 - _zz_when_ArraySlice_l113_383_4);
  assign _zz_when_ArraySlice_l113_383_1 = (_zz_when_ArraySlice_l113_383_2 + _zz_when_ArraySlice_l113_383_3);
  assign _zz_when_ArraySlice_l113_383_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_383_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_383_4 = {1'd0, _zz_when_ArraySlice_l112_383};
  assign _zz__zz_when_ArraySlice_l173_383 = (_zz__zz_when_ArraySlice_l173_383_1 + _zz__zz_when_ArraySlice_l173_383_2);
  assign _zz__zz_when_ArraySlice_l173_383_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_383_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_383_3 = {1'd0, _zz_when_ArraySlice_l112_383};
  assign _zz_when_ArraySlice_l118_383_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_383 = _zz_when_ArraySlice_l118_383_1[5:0];
  assign _zz_when_ArraySlice_l173_383_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_383_1 = {3'd0, _zz_when_ArraySlice_l173_383_2};
  assign _zz_when_ArraySlice_l173_383_3 = (_zz_when_ArraySlice_l173_383_4 + _zz_when_ArraySlice_l173_383_8);
  assign _zz_when_ArraySlice_l173_383_4 = (_zz_when_ArraySlice_l173_383 - _zz_when_ArraySlice_l173_383_5);
  assign _zz_when_ArraySlice_l173_383_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_383_7);
  assign _zz_when_ArraySlice_l173_383_5 = {1'd0, _zz_when_ArraySlice_l173_383_6};
  assign _zz_when_ArraySlice_l173_383_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_383_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l268_7_1 = (_zz_when_ArraySlice_l268_7_2 + _zz_when_ArraySlice_l268_7_7);
  assign _zz_when_ArraySlice_l268_7_2 = (_zz_when_ArraySlice_l268_7_3 + _zz_when_ArraySlice_l268_7_5);
  assign _zz_when_ArraySlice_l268_7_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l268_7_4);
  assign _zz_when_ArraySlice_l268_7_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l268_7_6 = 1'b1;
  assign _zz_when_ArraySlice_l268_7_5 = {5'd0, _zz_when_ArraySlice_l268_7_6};
  assign _zz_when_ArraySlice_l268_7_7 = (bReg * 3'b111);
  assign _zz_selectReadFifo_7_47 = 1'b1;
  assign _zz_selectReadFifo_7_46 = {5'd0, _zz_selectReadFifo_7_47};
  assign _zz_when_ArraySlice_l272_7 = (_zz_when_ArraySlice_l272_7_1 % aReg);
  assign _zz_when_ArraySlice_l272_7_1 = (handshakeTimes_7_value + _zz_when_ArraySlice_l272_7_2);
  assign _zz_when_ArraySlice_l272_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l272_7_2 = {12'd0, _zz_when_ArraySlice_l272_7_3};
  assign _zz_when_ArraySlice_l276_7_1 = (selectReadFifo_7 + _zz_when_ArraySlice_l276_7_2);
  assign _zz_when_ArraySlice_l276_7_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l277_7_1 = (_zz_when_ArraySlice_l277_7_2 - _zz_when_ArraySlice_l277_7_3);
  assign _zz_when_ArraySlice_l277_7 = {7'd0, _zz_when_ArraySlice_l277_7_1};
  assign _zz_when_ArraySlice_l277_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l277_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l277_7_3 = {5'd0, _zz_when_ArraySlice_l277_7_4};
  assign _zz__zz_when_ArraySlice_l94_46 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_46 = (_zz_when_ArraySlice_l95_46_1 - _zz_when_ArraySlice_l95_46_4);
  assign _zz_when_ArraySlice_l95_46_1 = (_zz_when_ArraySlice_l95_46_2 + _zz_when_ArraySlice_l95_46_3);
  assign _zz_when_ArraySlice_l95_46_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_46_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_46_4 = {1'd0, _zz_when_ArraySlice_l94_46};
  assign _zz__zz_when_ArraySlice_l279_7 = (_zz__zz_when_ArraySlice_l279_7_1 + _zz__zz_when_ArraySlice_l279_7_2);
  assign _zz__zz_when_ArraySlice_l279_7_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l279_7_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l279_7_3 = {1'd0, _zz_when_ArraySlice_l94_46};
  assign _zz_when_ArraySlice_l99_46_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_46 = _zz_when_ArraySlice_l99_46_1[5:0];
  assign _zz_when_ArraySlice_l279_7_1 = (outSliceNumb_7_value + _zz_when_ArraySlice_l279_7_2);
  assign _zz_when_ArraySlice_l279_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l279_7_2 = {6'd0, _zz_when_ArraySlice_l279_7_3};
  assign _zz_when_ArraySlice_l279_7_4 = (_zz_when_ArraySlice_l279_7 / aReg);
  assign _zz_selectReadFifo_7_48 = (selectReadFifo_7 - _zz_selectReadFifo_7_49);
  assign _zz_selectReadFifo_7_49 = {3'd0, bReg};
  assign _zz_selectReadFifo_7_51 = 1'b1;
  assign _zz_selectReadFifo_7_50 = {5'd0, _zz_selectReadFifo_7_51};
  assign _zz_selectReadFifo_7_52 = (selectReadFifo_7 + _zz_selectReadFifo_7_53);
  assign _zz_selectReadFifo_7_53 = (3'b111 * bReg);
  assign _zz_selectReadFifo_7_55 = 1'b1;
  assign _zz_selectReadFifo_7_54 = {5'd0, _zz_selectReadFifo_7_55};
  assign _zz_when_ArraySlice_l165_384 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_384_1);
  assign _zz_when_ArraySlice_l165_384_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_384_1 = {3'd0, _zz_when_ArraySlice_l165_384_2};
  assign _zz_when_ArraySlice_l166_384 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_384_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_384_3);
  assign _zz_when_ArraySlice_l166_384_1 = {1'd0, _zz_when_ArraySlice_l166_384_2};
  assign _zz_when_ArraySlice_l166_384_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_384_4);
  assign _zz_when_ArraySlice_l166_384_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_384_4 = {3'd0, _zz_when_ArraySlice_l166_384_5};
  assign _zz__zz_when_ArraySlice_l112_384 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_384 = (_zz_when_ArraySlice_l113_384_1 - _zz_when_ArraySlice_l113_384_4);
  assign _zz_when_ArraySlice_l113_384_1 = (_zz_when_ArraySlice_l113_384_2 + _zz_when_ArraySlice_l113_384_3);
  assign _zz_when_ArraySlice_l113_384_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_384_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_384_4 = {1'd0, _zz_when_ArraySlice_l112_384};
  assign _zz__zz_when_ArraySlice_l173_384 = (_zz__zz_when_ArraySlice_l173_384_1 + _zz__zz_when_ArraySlice_l173_384_2);
  assign _zz__zz_when_ArraySlice_l173_384_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_384_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_384_3 = {1'd0, _zz_when_ArraySlice_l112_384};
  assign _zz_when_ArraySlice_l118_384_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_384 = _zz_when_ArraySlice_l118_384_1[5:0];
  assign _zz_when_ArraySlice_l173_384_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_384_2 = (_zz_when_ArraySlice_l173_384_3 + _zz_when_ArraySlice_l173_384_8);
  assign _zz_when_ArraySlice_l173_384_3 = (_zz_when_ArraySlice_l173_384 - _zz_when_ArraySlice_l173_384_4);
  assign _zz_when_ArraySlice_l173_384_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_384_6);
  assign _zz_when_ArraySlice_l173_384_4 = {1'd0, _zz_when_ArraySlice_l173_384_5};
  assign _zz_when_ArraySlice_l173_384_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_384_6 = {3'd0, _zz_when_ArraySlice_l173_384_7};
  assign _zz_when_ArraySlice_l173_384_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_385 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_385_1);
  assign _zz_when_ArraySlice_l165_385_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_385_1 = {2'd0, _zz_when_ArraySlice_l165_385_2};
  assign _zz_when_ArraySlice_l166_385 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_385_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_385_2);
  assign _zz_when_ArraySlice_l166_385_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_385_3);
  assign _zz_when_ArraySlice_l166_385_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_385_3 = {2'd0, _zz_when_ArraySlice_l166_385_4};
  assign _zz__zz_when_ArraySlice_l112_385 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_385 = (_zz_when_ArraySlice_l113_385_1 - _zz_when_ArraySlice_l113_385_4);
  assign _zz_when_ArraySlice_l113_385_1 = (_zz_when_ArraySlice_l113_385_2 + _zz_when_ArraySlice_l113_385_3);
  assign _zz_when_ArraySlice_l113_385_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_385_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_385_4 = {1'd0, _zz_when_ArraySlice_l112_385};
  assign _zz__zz_when_ArraySlice_l173_385 = (_zz__zz_when_ArraySlice_l173_385_1 + _zz__zz_when_ArraySlice_l173_385_2);
  assign _zz__zz_when_ArraySlice_l173_385_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_385_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_385_3 = {1'd0, _zz_when_ArraySlice_l112_385};
  assign _zz_when_ArraySlice_l118_385_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_385 = _zz_when_ArraySlice_l118_385_1[5:0];
  assign _zz_when_ArraySlice_l173_385_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_385_1 = {1'd0, _zz_when_ArraySlice_l173_385_2};
  assign _zz_when_ArraySlice_l173_385_3 = (_zz_when_ArraySlice_l173_385_4 + _zz_when_ArraySlice_l173_385_9);
  assign _zz_when_ArraySlice_l173_385_4 = (_zz_when_ArraySlice_l173_385 - _zz_when_ArraySlice_l173_385_5);
  assign _zz_when_ArraySlice_l173_385_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_385_7);
  assign _zz_when_ArraySlice_l173_385_5 = {1'd0, _zz_when_ArraySlice_l173_385_6};
  assign _zz_when_ArraySlice_l173_385_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_385_7 = {2'd0, _zz_when_ArraySlice_l173_385_8};
  assign _zz_when_ArraySlice_l173_385_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_386 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_386_1);
  assign _zz_when_ArraySlice_l165_386_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_386_1 = {1'd0, _zz_when_ArraySlice_l165_386_2};
  assign _zz_when_ArraySlice_l166_386 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_386_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_386_2);
  assign _zz_when_ArraySlice_l166_386_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_386_3);
  assign _zz_when_ArraySlice_l166_386_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_386_3 = {1'd0, _zz_when_ArraySlice_l166_386_4};
  assign _zz__zz_when_ArraySlice_l112_386 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_386 = (_zz_when_ArraySlice_l113_386_1 - _zz_when_ArraySlice_l113_386_4);
  assign _zz_when_ArraySlice_l113_386_1 = (_zz_when_ArraySlice_l113_386_2 + _zz_when_ArraySlice_l113_386_3);
  assign _zz_when_ArraySlice_l113_386_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_386_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_386_4 = {1'd0, _zz_when_ArraySlice_l112_386};
  assign _zz__zz_when_ArraySlice_l173_386 = (_zz__zz_when_ArraySlice_l173_386_1 + _zz__zz_when_ArraySlice_l173_386_2);
  assign _zz__zz_when_ArraySlice_l173_386_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_386_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_386_3 = {1'd0, _zz_when_ArraySlice_l112_386};
  assign _zz_when_ArraySlice_l118_386_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_386 = _zz_when_ArraySlice_l118_386_1[5:0];
  assign _zz_when_ArraySlice_l173_386_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_386_1 = {1'd0, _zz_when_ArraySlice_l173_386_2};
  assign _zz_when_ArraySlice_l173_386_3 = (_zz_when_ArraySlice_l173_386_4 + _zz_when_ArraySlice_l173_386_9);
  assign _zz_when_ArraySlice_l173_386_4 = (_zz_when_ArraySlice_l173_386 - _zz_when_ArraySlice_l173_386_5);
  assign _zz_when_ArraySlice_l173_386_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_386_7);
  assign _zz_when_ArraySlice_l173_386_5 = {1'd0, _zz_when_ArraySlice_l173_386_6};
  assign _zz_when_ArraySlice_l173_386_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_386_7 = {1'd0, _zz_when_ArraySlice_l173_386_8};
  assign _zz_when_ArraySlice_l173_386_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_387 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_387_1);
  assign _zz_when_ArraySlice_l165_387_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_387_1 = {1'd0, _zz_when_ArraySlice_l165_387_2};
  assign _zz_when_ArraySlice_l166_387 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_387_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_387_2);
  assign _zz_when_ArraySlice_l166_387_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_387_3);
  assign _zz_when_ArraySlice_l166_387_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_387_3 = {1'd0, _zz_when_ArraySlice_l166_387_4};
  assign _zz__zz_when_ArraySlice_l112_387 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_387 = (_zz_when_ArraySlice_l113_387_1 - _zz_when_ArraySlice_l113_387_4);
  assign _zz_when_ArraySlice_l113_387_1 = (_zz_when_ArraySlice_l113_387_2 + _zz_when_ArraySlice_l113_387_3);
  assign _zz_when_ArraySlice_l113_387_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_387_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_387_4 = {1'd0, _zz_when_ArraySlice_l112_387};
  assign _zz__zz_when_ArraySlice_l173_387 = (_zz__zz_when_ArraySlice_l173_387_1 + _zz__zz_when_ArraySlice_l173_387_2);
  assign _zz__zz_when_ArraySlice_l173_387_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_387_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_387_3 = {1'd0, _zz_when_ArraySlice_l112_387};
  assign _zz_when_ArraySlice_l118_387_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_387 = _zz_when_ArraySlice_l118_387_1[5:0];
  assign _zz_when_ArraySlice_l173_387_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_387_1 = {1'd0, _zz_when_ArraySlice_l173_387_2};
  assign _zz_when_ArraySlice_l173_387_3 = (_zz_when_ArraySlice_l173_387_4 + _zz_when_ArraySlice_l173_387_9);
  assign _zz_when_ArraySlice_l173_387_4 = (_zz_when_ArraySlice_l173_387 - _zz_when_ArraySlice_l173_387_5);
  assign _zz_when_ArraySlice_l173_387_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_387_7);
  assign _zz_when_ArraySlice_l173_387_5 = {1'd0, _zz_when_ArraySlice_l173_387_6};
  assign _zz_when_ArraySlice_l173_387_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_387_7 = {1'd0, _zz_when_ArraySlice_l173_387_8};
  assign _zz_when_ArraySlice_l173_387_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_388 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_388_1);
  assign _zz_when_ArraySlice_l165_388_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_388 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_388_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_388_2);
  assign _zz_when_ArraySlice_l166_388_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_388_3);
  assign _zz_when_ArraySlice_l166_388_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_388 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_388 = (_zz_when_ArraySlice_l113_388_1 - _zz_when_ArraySlice_l113_388_4);
  assign _zz_when_ArraySlice_l113_388_1 = (_zz_when_ArraySlice_l113_388_2 + _zz_when_ArraySlice_l113_388_3);
  assign _zz_when_ArraySlice_l113_388_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_388_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_388_4 = {1'd0, _zz_when_ArraySlice_l112_388};
  assign _zz__zz_when_ArraySlice_l173_388 = (_zz__zz_when_ArraySlice_l173_388_1 + _zz__zz_when_ArraySlice_l173_388_2);
  assign _zz__zz_when_ArraySlice_l173_388_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_388_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_388_3 = {1'd0, _zz_when_ArraySlice_l112_388};
  assign _zz_when_ArraySlice_l118_388_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_388 = _zz_when_ArraySlice_l118_388_1[5:0];
  assign _zz_when_ArraySlice_l173_388_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_388_1 = {1'd0, _zz_when_ArraySlice_l173_388_2};
  assign _zz_when_ArraySlice_l173_388_3 = (_zz_when_ArraySlice_l173_388_4 + _zz_when_ArraySlice_l173_388_8);
  assign _zz_when_ArraySlice_l173_388_4 = (_zz_when_ArraySlice_l173_388 - _zz_when_ArraySlice_l173_388_5);
  assign _zz_when_ArraySlice_l173_388_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_388_7);
  assign _zz_when_ArraySlice_l173_388_5 = {1'd0, _zz_when_ArraySlice_l173_388_6};
  assign _zz_when_ArraySlice_l173_388_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_388_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_389 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_389_1);
  assign _zz_when_ArraySlice_l165_389_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_389_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_389 = {1'd0, _zz_when_ArraySlice_l166_389_1};
  assign _zz_when_ArraySlice_l166_389_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_389_3);
  assign _zz_when_ArraySlice_l166_389_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_389_4);
  assign _zz_when_ArraySlice_l166_389_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_389 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_389 = (_zz_when_ArraySlice_l113_389_1 - _zz_when_ArraySlice_l113_389_4);
  assign _zz_when_ArraySlice_l113_389_1 = (_zz_when_ArraySlice_l113_389_2 + _zz_when_ArraySlice_l113_389_3);
  assign _zz_when_ArraySlice_l113_389_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_389_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_389_4 = {1'd0, _zz_when_ArraySlice_l112_389};
  assign _zz__zz_when_ArraySlice_l173_389 = (_zz__zz_when_ArraySlice_l173_389_1 + _zz__zz_when_ArraySlice_l173_389_2);
  assign _zz__zz_when_ArraySlice_l173_389_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_389_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_389_3 = {1'd0, _zz_when_ArraySlice_l112_389};
  assign _zz_when_ArraySlice_l118_389_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_389 = _zz_when_ArraySlice_l118_389_1[5:0];
  assign _zz_when_ArraySlice_l173_389_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_389_1 = {2'd0, _zz_when_ArraySlice_l173_389_2};
  assign _zz_when_ArraySlice_l173_389_3 = (_zz_when_ArraySlice_l173_389_4 + _zz_when_ArraySlice_l173_389_8);
  assign _zz_when_ArraySlice_l173_389_4 = (_zz_when_ArraySlice_l173_389 - _zz_when_ArraySlice_l173_389_5);
  assign _zz_when_ArraySlice_l173_389_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_389_7);
  assign _zz_when_ArraySlice_l173_389_5 = {1'd0, _zz_when_ArraySlice_l173_389_6};
  assign _zz_when_ArraySlice_l173_389_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_389_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_390 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_390_1);
  assign _zz_when_ArraySlice_l165_390_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_390_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_390 = {1'd0, _zz_when_ArraySlice_l166_390_1};
  assign _zz_when_ArraySlice_l166_390_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_390_3);
  assign _zz_when_ArraySlice_l166_390_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_390_4);
  assign _zz_when_ArraySlice_l166_390_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_390 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_390 = (_zz_when_ArraySlice_l113_390_1 - _zz_when_ArraySlice_l113_390_4);
  assign _zz_when_ArraySlice_l113_390_1 = (_zz_when_ArraySlice_l113_390_2 + _zz_when_ArraySlice_l113_390_3);
  assign _zz_when_ArraySlice_l113_390_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_390_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_390_4 = {1'd0, _zz_when_ArraySlice_l112_390};
  assign _zz__zz_when_ArraySlice_l173_390 = (_zz__zz_when_ArraySlice_l173_390_1 + _zz__zz_when_ArraySlice_l173_390_2);
  assign _zz__zz_when_ArraySlice_l173_390_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_390_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_390_3 = {1'd0, _zz_when_ArraySlice_l112_390};
  assign _zz_when_ArraySlice_l118_390_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_390 = _zz_when_ArraySlice_l118_390_1[5:0];
  assign _zz_when_ArraySlice_l173_390_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_390_1 = {2'd0, _zz_when_ArraySlice_l173_390_2};
  assign _zz_when_ArraySlice_l173_390_3 = (_zz_when_ArraySlice_l173_390_4 + _zz_when_ArraySlice_l173_390_8);
  assign _zz_when_ArraySlice_l173_390_4 = (_zz_when_ArraySlice_l173_390 - _zz_when_ArraySlice_l173_390_5);
  assign _zz_when_ArraySlice_l173_390_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_390_7);
  assign _zz_when_ArraySlice_l173_390_5 = {1'd0, _zz_when_ArraySlice_l173_390_6};
  assign _zz_when_ArraySlice_l173_390_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_390_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_391 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_391_1);
  assign _zz_when_ArraySlice_l165_391_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_391_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_391 = {2'd0, _zz_when_ArraySlice_l166_391_1};
  assign _zz_when_ArraySlice_l166_391_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_391_3);
  assign _zz_when_ArraySlice_l166_391_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_391_4);
  assign _zz_when_ArraySlice_l166_391_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_391 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_391 = (_zz_when_ArraySlice_l113_391_1 - _zz_when_ArraySlice_l113_391_4);
  assign _zz_when_ArraySlice_l113_391_1 = (_zz_when_ArraySlice_l113_391_2 + _zz_when_ArraySlice_l113_391_3);
  assign _zz_when_ArraySlice_l113_391_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_391_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_391_4 = {1'd0, _zz_when_ArraySlice_l112_391};
  assign _zz__zz_when_ArraySlice_l173_391 = (_zz__zz_when_ArraySlice_l173_391_1 + _zz__zz_when_ArraySlice_l173_391_2);
  assign _zz__zz_when_ArraySlice_l173_391_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_391_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_391_3 = {1'd0, _zz_when_ArraySlice_l112_391};
  assign _zz_when_ArraySlice_l118_391_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_391 = _zz_when_ArraySlice_l118_391_1[5:0];
  assign _zz_when_ArraySlice_l173_391_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_391_1 = {3'd0, _zz_when_ArraySlice_l173_391_2};
  assign _zz_when_ArraySlice_l173_391_3 = (_zz_when_ArraySlice_l173_391_4 + _zz_when_ArraySlice_l173_391_8);
  assign _zz_when_ArraySlice_l173_391_4 = (_zz_when_ArraySlice_l173_391 - _zz_when_ArraySlice_l173_391_5);
  assign _zz_when_ArraySlice_l173_391_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_391_7);
  assign _zz_when_ArraySlice_l173_391_5 = {1'd0, _zz_when_ArraySlice_l173_391_6};
  assign _zz_when_ArraySlice_l173_391_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_391_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l288_7_1 = (_zz_when_ArraySlice_l288_7_2 + _zz_when_ArraySlice_l288_7_7);
  assign _zz_when_ArraySlice_l288_7_2 = (_zz_when_ArraySlice_l288_7_3 + _zz_when_ArraySlice_l288_7_5);
  assign _zz_when_ArraySlice_l288_7_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l288_7_4);
  assign _zz_when_ArraySlice_l288_7_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_7_6 = 1'b1;
  assign _zz_when_ArraySlice_l288_7_5 = {5'd0, _zz_when_ArraySlice_l288_7_6};
  assign _zz_when_ArraySlice_l288_7_7 = (bReg * 3'b111);
  assign _zz_selectReadFifo_7_57 = 1'b1;
  assign _zz_selectReadFifo_7_56 = {5'd0, _zz_selectReadFifo_7_57};
  assign _zz_when_ArraySlice_l292_7 = (_zz_when_ArraySlice_l292_7_1 % aReg);
  assign _zz_when_ArraySlice_l292_7_1 = (handshakeTimes_7_value + _zz_when_ArraySlice_l292_7_2);
  assign _zz_when_ArraySlice_l292_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l292_7_2 = {12'd0, _zz_when_ArraySlice_l292_7_3};
  assign _zz_when_ArraySlice_l303_7_1 = (_zz_when_ArraySlice_l303_7_2 - _zz_when_ArraySlice_l303_7_3);
  assign _zz_when_ArraySlice_l303_7 = {7'd0, _zz_when_ArraySlice_l303_7_1};
  assign _zz_when_ArraySlice_l303_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l303_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l303_7_3 = {5'd0, _zz_when_ArraySlice_l303_7_4};
  assign _zz__zz_when_ArraySlice_l94_47 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_47 = (_zz_when_ArraySlice_l95_47_1 - _zz_when_ArraySlice_l95_47_4);
  assign _zz_when_ArraySlice_l95_47_1 = (_zz_when_ArraySlice_l95_47_2 + _zz_when_ArraySlice_l95_47_3);
  assign _zz_when_ArraySlice_l95_47_2 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l95_47_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l95_47_4 = {1'd0, _zz_when_ArraySlice_l94_47};
  assign _zz__zz_when_ArraySlice_l304_7 = (_zz__zz_when_ArraySlice_l304_7_1 + _zz__zz_when_ArraySlice_l304_7_2);
  assign _zz__zz_when_ArraySlice_l304_7_1 = {1'd0, hReg};
  assign _zz__zz_when_ArraySlice_l304_7_2 = (aReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l304_7_3 = {1'd0, _zz_when_ArraySlice_l94_47};
  assign _zz_when_ArraySlice_l99_47_1 = 7'h40;
  assign _zz_when_ArraySlice_l99_47 = _zz_when_ArraySlice_l99_47_1[5:0];
  assign _zz_when_ArraySlice_l304_7_1 = (outSliceNumb_7_value + _zz_when_ArraySlice_l304_7_2);
  assign _zz_when_ArraySlice_l304_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l304_7_2 = {6'd0, _zz_when_ArraySlice_l304_7_3};
  assign _zz_when_ArraySlice_l304_7_4 = (_zz_when_ArraySlice_l304_7 / aReg);
  assign _zz_selectReadFifo_7_58 = (selectReadFifo_7 - _zz_selectReadFifo_7_59);
  assign _zz_selectReadFifo_7_59 = {3'd0, bReg};
  assign _zz_selectReadFifo_7_61 = 1'b1;
  assign _zz_selectReadFifo_7_60 = {5'd0, _zz_selectReadFifo_7_61};
  assign _zz_when_ArraySlice_l165_392 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_392_1);
  assign _zz_when_ArraySlice_l165_392_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_392_1 = {3'd0, _zz_when_ArraySlice_l165_392_2};
  assign _zz_when_ArraySlice_l166_392 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_392_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_392_3);
  assign _zz_when_ArraySlice_l166_392_1 = {1'd0, _zz_when_ArraySlice_l166_392_2};
  assign _zz_when_ArraySlice_l166_392_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_392_4);
  assign _zz_when_ArraySlice_l166_392_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_392_4 = {3'd0, _zz_when_ArraySlice_l166_392_5};
  assign _zz__zz_when_ArraySlice_l112_392 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_392 = (_zz_when_ArraySlice_l113_392_1 - _zz_when_ArraySlice_l113_392_4);
  assign _zz_when_ArraySlice_l113_392_1 = (_zz_when_ArraySlice_l113_392_2 + _zz_when_ArraySlice_l113_392_3);
  assign _zz_when_ArraySlice_l113_392_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_392_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_392_4 = {1'd0, _zz_when_ArraySlice_l112_392};
  assign _zz__zz_when_ArraySlice_l173_392 = (_zz__zz_when_ArraySlice_l173_392_1 + _zz__zz_when_ArraySlice_l173_392_2);
  assign _zz__zz_when_ArraySlice_l173_392_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_392_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_392_3 = {1'd0, _zz_when_ArraySlice_l112_392};
  assign _zz_when_ArraySlice_l118_392_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_392 = _zz_when_ArraySlice_l118_392_1[5:0];
  assign _zz_when_ArraySlice_l173_392_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_392_2 = (_zz_when_ArraySlice_l173_392_3 + _zz_when_ArraySlice_l173_392_8);
  assign _zz_when_ArraySlice_l173_392_3 = (_zz_when_ArraySlice_l173_392 - _zz_when_ArraySlice_l173_392_4);
  assign _zz_when_ArraySlice_l173_392_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_392_6);
  assign _zz_when_ArraySlice_l173_392_4 = {1'd0, _zz_when_ArraySlice_l173_392_5};
  assign _zz_when_ArraySlice_l173_392_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_392_6 = {3'd0, _zz_when_ArraySlice_l173_392_7};
  assign _zz_when_ArraySlice_l173_392_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_393 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_393_1);
  assign _zz_when_ArraySlice_l165_393_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_393_1 = {2'd0, _zz_when_ArraySlice_l165_393_2};
  assign _zz_when_ArraySlice_l166_393 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_393_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_393_2);
  assign _zz_when_ArraySlice_l166_393_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_393_3);
  assign _zz_when_ArraySlice_l166_393_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_393_3 = {2'd0, _zz_when_ArraySlice_l166_393_4};
  assign _zz__zz_when_ArraySlice_l112_393 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_393 = (_zz_when_ArraySlice_l113_393_1 - _zz_when_ArraySlice_l113_393_4);
  assign _zz_when_ArraySlice_l113_393_1 = (_zz_when_ArraySlice_l113_393_2 + _zz_when_ArraySlice_l113_393_3);
  assign _zz_when_ArraySlice_l113_393_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_393_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_393_4 = {1'd0, _zz_when_ArraySlice_l112_393};
  assign _zz__zz_when_ArraySlice_l173_393 = (_zz__zz_when_ArraySlice_l173_393_1 + _zz__zz_when_ArraySlice_l173_393_2);
  assign _zz__zz_when_ArraySlice_l173_393_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_393_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_393_3 = {1'd0, _zz_when_ArraySlice_l112_393};
  assign _zz_when_ArraySlice_l118_393_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_393 = _zz_when_ArraySlice_l118_393_1[5:0];
  assign _zz_when_ArraySlice_l173_393_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_393_1 = {1'd0, _zz_when_ArraySlice_l173_393_2};
  assign _zz_when_ArraySlice_l173_393_3 = (_zz_when_ArraySlice_l173_393_4 + _zz_when_ArraySlice_l173_393_9);
  assign _zz_when_ArraySlice_l173_393_4 = (_zz_when_ArraySlice_l173_393 - _zz_when_ArraySlice_l173_393_5);
  assign _zz_when_ArraySlice_l173_393_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_393_7);
  assign _zz_when_ArraySlice_l173_393_5 = {1'd0, _zz_when_ArraySlice_l173_393_6};
  assign _zz_when_ArraySlice_l173_393_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_393_7 = {2'd0, _zz_when_ArraySlice_l173_393_8};
  assign _zz_when_ArraySlice_l173_393_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_394 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_394_1);
  assign _zz_when_ArraySlice_l165_394_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_394_1 = {1'd0, _zz_when_ArraySlice_l165_394_2};
  assign _zz_when_ArraySlice_l166_394 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_394_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_394_2);
  assign _zz_when_ArraySlice_l166_394_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_394_3);
  assign _zz_when_ArraySlice_l166_394_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_394_3 = {1'd0, _zz_when_ArraySlice_l166_394_4};
  assign _zz__zz_when_ArraySlice_l112_394 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_394 = (_zz_when_ArraySlice_l113_394_1 - _zz_when_ArraySlice_l113_394_4);
  assign _zz_when_ArraySlice_l113_394_1 = (_zz_when_ArraySlice_l113_394_2 + _zz_when_ArraySlice_l113_394_3);
  assign _zz_when_ArraySlice_l113_394_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_394_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_394_4 = {1'd0, _zz_when_ArraySlice_l112_394};
  assign _zz__zz_when_ArraySlice_l173_394 = (_zz__zz_when_ArraySlice_l173_394_1 + _zz__zz_when_ArraySlice_l173_394_2);
  assign _zz__zz_when_ArraySlice_l173_394_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_394_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_394_3 = {1'd0, _zz_when_ArraySlice_l112_394};
  assign _zz_when_ArraySlice_l118_394_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_394 = _zz_when_ArraySlice_l118_394_1[5:0];
  assign _zz_when_ArraySlice_l173_394_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_394_1 = {1'd0, _zz_when_ArraySlice_l173_394_2};
  assign _zz_when_ArraySlice_l173_394_3 = (_zz_when_ArraySlice_l173_394_4 + _zz_when_ArraySlice_l173_394_9);
  assign _zz_when_ArraySlice_l173_394_4 = (_zz_when_ArraySlice_l173_394 - _zz_when_ArraySlice_l173_394_5);
  assign _zz_when_ArraySlice_l173_394_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_394_7);
  assign _zz_when_ArraySlice_l173_394_5 = {1'd0, _zz_when_ArraySlice_l173_394_6};
  assign _zz_when_ArraySlice_l173_394_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_394_7 = {1'd0, _zz_when_ArraySlice_l173_394_8};
  assign _zz_when_ArraySlice_l173_394_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_395 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_395_1);
  assign _zz_when_ArraySlice_l165_395_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_395_1 = {1'd0, _zz_when_ArraySlice_l165_395_2};
  assign _zz_when_ArraySlice_l166_395 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_395_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_395_2);
  assign _zz_when_ArraySlice_l166_395_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_395_3);
  assign _zz_when_ArraySlice_l166_395_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_395_3 = {1'd0, _zz_when_ArraySlice_l166_395_4};
  assign _zz__zz_when_ArraySlice_l112_395 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_395 = (_zz_when_ArraySlice_l113_395_1 - _zz_when_ArraySlice_l113_395_4);
  assign _zz_when_ArraySlice_l113_395_1 = (_zz_when_ArraySlice_l113_395_2 + _zz_when_ArraySlice_l113_395_3);
  assign _zz_when_ArraySlice_l113_395_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_395_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_395_4 = {1'd0, _zz_when_ArraySlice_l112_395};
  assign _zz__zz_when_ArraySlice_l173_395 = (_zz__zz_when_ArraySlice_l173_395_1 + _zz__zz_when_ArraySlice_l173_395_2);
  assign _zz__zz_when_ArraySlice_l173_395_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_395_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_395_3 = {1'd0, _zz_when_ArraySlice_l112_395};
  assign _zz_when_ArraySlice_l118_395_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_395 = _zz_when_ArraySlice_l118_395_1[5:0];
  assign _zz_when_ArraySlice_l173_395_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_395_1 = {1'd0, _zz_when_ArraySlice_l173_395_2};
  assign _zz_when_ArraySlice_l173_395_3 = (_zz_when_ArraySlice_l173_395_4 + _zz_when_ArraySlice_l173_395_9);
  assign _zz_when_ArraySlice_l173_395_4 = (_zz_when_ArraySlice_l173_395 - _zz_when_ArraySlice_l173_395_5);
  assign _zz_when_ArraySlice_l173_395_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_395_7);
  assign _zz_when_ArraySlice_l173_395_5 = {1'd0, _zz_when_ArraySlice_l173_395_6};
  assign _zz_when_ArraySlice_l173_395_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_395_7 = {1'd0, _zz_when_ArraySlice_l173_395_8};
  assign _zz_when_ArraySlice_l173_395_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_396 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_396_1);
  assign _zz_when_ArraySlice_l165_396_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_396 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_396_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_396_2);
  assign _zz_when_ArraySlice_l166_396_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_396_3);
  assign _zz_when_ArraySlice_l166_396_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_396 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_396 = (_zz_when_ArraySlice_l113_396_1 - _zz_when_ArraySlice_l113_396_4);
  assign _zz_when_ArraySlice_l113_396_1 = (_zz_when_ArraySlice_l113_396_2 + _zz_when_ArraySlice_l113_396_3);
  assign _zz_when_ArraySlice_l113_396_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_396_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_396_4 = {1'd0, _zz_when_ArraySlice_l112_396};
  assign _zz__zz_when_ArraySlice_l173_396 = (_zz__zz_when_ArraySlice_l173_396_1 + _zz__zz_when_ArraySlice_l173_396_2);
  assign _zz__zz_when_ArraySlice_l173_396_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_396_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_396_3 = {1'd0, _zz_when_ArraySlice_l112_396};
  assign _zz_when_ArraySlice_l118_396_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_396 = _zz_when_ArraySlice_l118_396_1[5:0];
  assign _zz_when_ArraySlice_l173_396_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_396_1 = {1'd0, _zz_when_ArraySlice_l173_396_2};
  assign _zz_when_ArraySlice_l173_396_3 = (_zz_when_ArraySlice_l173_396_4 + _zz_when_ArraySlice_l173_396_8);
  assign _zz_when_ArraySlice_l173_396_4 = (_zz_when_ArraySlice_l173_396 - _zz_when_ArraySlice_l173_396_5);
  assign _zz_when_ArraySlice_l173_396_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_396_7);
  assign _zz_when_ArraySlice_l173_396_5 = {1'd0, _zz_when_ArraySlice_l173_396_6};
  assign _zz_when_ArraySlice_l173_396_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_396_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_397 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_397_1);
  assign _zz_when_ArraySlice_l165_397_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_397_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_397 = {1'd0, _zz_when_ArraySlice_l166_397_1};
  assign _zz_when_ArraySlice_l166_397_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_397_3);
  assign _zz_when_ArraySlice_l166_397_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_397_4);
  assign _zz_when_ArraySlice_l166_397_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_397 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_397 = (_zz_when_ArraySlice_l113_397_1 - _zz_when_ArraySlice_l113_397_4);
  assign _zz_when_ArraySlice_l113_397_1 = (_zz_when_ArraySlice_l113_397_2 + _zz_when_ArraySlice_l113_397_3);
  assign _zz_when_ArraySlice_l113_397_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_397_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_397_4 = {1'd0, _zz_when_ArraySlice_l112_397};
  assign _zz__zz_when_ArraySlice_l173_397 = (_zz__zz_when_ArraySlice_l173_397_1 + _zz__zz_when_ArraySlice_l173_397_2);
  assign _zz__zz_when_ArraySlice_l173_397_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_397_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_397_3 = {1'd0, _zz_when_ArraySlice_l112_397};
  assign _zz_when_ArraySlice_l118_397_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_397 = _zz_when_ArraySlice_l118_397_1[5:0];
  assign _zz_when_ArraySlice_l173_397_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_397_1 = {2'd0, _zz_when_ArraySlice_l173_397_2};
  assign _zz_when_ArraySlice_l173_397_3 = (_zz_when_ArraySlice_l173_397_4 + _zz_when_ArraySlice_l173_397_8);
  assign _zz_when_ArraySlice_l173_397_4 = (_zz_when_ArraySlice_l173_397 - _zz_when_ArraySlice_l173_397_5);
  assign _zz_when_ArraySlice_l173_397_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_397_7);
  assign _zz_when_ArraySlice_l173_397_5 = {1'd0, _zz_when_ArraySlice_l173_397_6};
  assign _zz_when_ArraySlice_l173_397_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_397_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_398 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_398_1);
  assign _zz_when_ArraySlice_l165_398_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_398_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_398 = {1'd0, _zz_when_ArraySlice_l166_398_1};
  assign _zz_when_ArraySlice_l166_398_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_398_3);
  assign _zz_when_ArraySlice_l166_398_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_398_4);
  assign _zz_when_ArraySlice_l166_398_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_398 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_398 = (_zz_when_ArraySlice_l113_398_1 - _zz_when_ArraySlice_l113_398_4);
  assign _zz_when_ArraySlice_l113_398_1 = (_zz_when_ArraySlice_l113_398_2 + _zz_when_ArraySlice_l113_398_3);
  assign _zz_when_ArraySlice_l113_398_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_398_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_398_4 = {1'd0, _zz_when_ArraySlice_l112_398};
  assign _zz__zz_when_ArraySlice_l173_398 = (_zz__zz_when_ArraySlice_l173_398_1 + _zz__zz_when_ArraySlice_l173_398_2);
  assign _zz__zz_when_ArraySlice_l173_398_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_398_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_398_3 = {1'd0, _zz_when_ArraySlice_l112_398};
  assign _zz_when_ArraySlice_l118_398_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_398 = _zz_when_ArraySlice_l118_398_1[5:0];
  assign _zz_when_ArraySlice_l173_398_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_398_1 = {2'd0, _zz_when_ArraySlice_l173_398_2};
  assign _zz_when_ArraySlice_l173_398_3 = (_zz_when_ArraySlice_l173_398_4 + _zz_when_ArraySlice_l173_398_8);
  assign _zz_when_ArraySlice_l173_398_4 = (_zz_when_ArraySlice_l173_398 - _zz_when_ArraySlice_l173_398_5);
  assign _zz_when_ArraySlice_l173_398_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_398_7);
  assign _zz_when_ArraySlice_l173_398_5 = {1'd0, _zz_when_ArraySlice_l173_398_6};
  assign _zz_when_ArraySlice_l173_398_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_398_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_399 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_399_1);
  assign _zz_when_ArraySlice_l165_399_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_399_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_399 = {2'd0, _zz_when_ArraySlice_l166_399_1};
  assign _zz_when_ArraySlice_l166_399_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_399_3);
  assign _zz_when_ArraySlice_l166_399_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_399_4);
  assign _zz_when_ArraySlice_l166_399_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_399 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_399 = (_zz_when_ArraySlice_l113_399_1 - _zz_when_ArraySlice_l113_399_4);
  assign _zz_when_ArraySlice_l113_399_1 = (_zz_when_ArraySlice_l113_399_2 + _zz_when_ArraySlice_l113_399_3);
  assign _zz_when_ArraySlice_l113_399_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_399_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_399_4 = {1'd0, _zz_when_ArraySlice_l112_399};
  assign _zz__zz_when_ArraySlice_l173_399 = (_zz__zz_when_ArraySlice_l173_399_1 + _zz__zz_when_ArraySlice_l173_399_2);
  assign _zz__zz_when_ArraySlice_l173_399_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_399_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_399_3 = {1'd0, _zz_when_ArraySlice_l112_399};
  assign _zz_when_ArraySlice_l118_399_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_399 = _zz_when_ArraySlice_l118_399_1[5:0];
  assign _zz_when_ArraySlice_l173_399_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_399_1 = {3'd0, _zz_when_ArraySlice_l173_399_2};
  assign _zz_when_ArraySlice_l173_399_3 = (_zz_when_ArraySlice_l173_399_4 + _zz_when_ArraySlice_l173_399_8);
  assign _zz_when_ArraySlice_l173_399_4 = (_zz_when_ArraySlice_l173_399 - _zz_when_ArraySlice_l173_399_5);
  assign _zz_when_ArraySlice_l173_399_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_399_7);
  assign _zz_when_ArraySlice_l173_399_5 = {1'd0, _zz_when_ArraySlice_l173_399_6};
  assign _zz_when_ArraySlice_l173_399_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_399_8 = {1'd0, selectWriteFifo};
  assign _zz_selectReadFifo_7_63 = 1'b1;
  assign _zz_selectReadFifo_7_62 = {5'd0, _zz_selectReadFifo_7_63};
  assign _zz_when_ArraySlice_l315_7 = (_zz_when_ArraySlice_l315_7_1 % aReg);
  assign _zz_when_ArraySlice_l315_7_1 = (handshakeTimes_7_value + _zz_when_ArraySlice_l315_7_2);
  assign _zz_when_ArraySlice_l315_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l315_7_2 = {12'd0, _zz_when_ArraySlice_l315_7_3};
  assign _zz_when_ArraySlice_l301_7 = (selectReadFifo_7 + _zz_when_ArraySlice_l301_7_1);
  assign _zz_when_ArraySlice_l301_7_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l322_7_1 = (_zz_when_ArraySlice_l322_7_2 - _zz_when_ArraySlice_l322_7_3);
  assign _zz_when_ArraySlice_l322_7 = {7'd0, _zz_when_ArraySlice_l322_7_1};
  assign _zz_when_ArraySlice_l322_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l322_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l322_7_3 = {5'd0, _zz_when_ArraySlice_l322_7_4};
  assign _zz_when_ArraySlice_l189 = (selectReadFifo_0 - _zz_when_ArraySlice_l189_1);
  assign _zz_when_ArraySlice_l189_1 = (selectReadFifo_0 % bReg);
  assign _zz_when_ArraySlice_l189_1_1 = (selectReadFifo_1 - _zz_when_ArraySlice_l189_1_2);
  assign _zz_when_ArraySlice_l189_1_2 = (selectReadFifo_1 % bReg);
  assign _zz_when_ArraySlice_l189_2 = (selectReadFifo_2 - _zz_when_ArraySlice_l189_2_1);
  assign _zz_when_ArraySlice_l189_2_1 = (selectReadFifo_2 % bReg);
  assign _zz_when_ArraySlice_l189_3 = (selectReadFifo_3 - _zz_when_ArraySlice_l189_3_1);
  assign _zz_when_ArraySlice_l189_3_1 = (selectReadFifo_3 % bReg);
  assign _zz_when_ArraySlice_l189_4 = (selectReadFifo_4 - _zz_when_ArraySlice_l189_4_1);
  assign _zz_when_ArraySlice_l189_4_1 = (selectReadFifo_4 % bReg);
  assign _zz_when_ArraySlice_l189_5 = (selectReadFifo_5 - _zz_when_ArraySlice_l189_5_1);
  assign _zz_when_ArraySlice_l189_5_1 = (selectReadFifo_5 % bReg);
  assign _zz_when_ArraySlice_l189_6 = (selectReadFifo_6 - _zz_when_ArraySlice_l189_6_1);
  assign _zz_when_ArraySlice_l189_6_1 = (selectReadFifo_6 % bReg);
  assign _zz_when_ArraySlice_l189_7 = (selectReadFifo_7 - _zz_when_ArraySlice_l189_7_1);
  assign _zz_when_ArraySlice_l189_7_1 = (selectReadFifo_7 % bReg);
  assign _zz_when_ArraySlice_l334_1 = {1'd0, hReg};
  assign _zz_when_ArraySlice_l338_2 = (hReg - _zz_when_ArraySlice_l338_3);
  assign _zz_when_ArraySlice_l338_1 = {1'd0, _zz_when_ArraySlice_l338_2};
  assign _zz_when_ArraySlice_l338_4 = 1'b1;
  assign _zz_when_ArraySlice_l338_3 = {5'd0, _zz_when_ArraySlice_l338_4};
  assign _zz_when_ArraySlice_l339 = (wReg - _zz_when_ArraySlice_l339_1);
  assign _zz_when_ArraySlice_l339_2 = 1'b1;
  assign _zz_when_ArraySlice_l339_1 = {5'd0, _zz_when_ArraySlice_l339_2};
  assign _zz_selectWriteFifo_3 = 1'b1;
  assign _zz_selectWriteFifo_2 = {5'd0, _zz_selectWriteFifo_3};
  assign _zz_when_ArraySlice_l165_400 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_400_1);
  assign _zz_when_ArraySlice_l165_400_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_400_1 = {3'd0, _zz_when_ArraySlice_l165_400_2};
  assign _zz_when_ArraySlice_l166_400 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_400_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_400_3);
  assign _zz_when_ArraySlice_l166_400_1 = {1'd0, _zz_when_ArraySlice_l166_400_2};
  assign _zz_when_ArraySlice_l166_400_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_400_4);
  assign _zz_when_ArraySlice_l166_400_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_400_4 = {3'd0, _zz_when_ArraySlice_l166_400_5};
  assign _zz__zz_when_ArraySlice_l112_400 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_400 = (_zz_when_ArraySlice_l113_400_1 - _zz_when_ArraySlice_l113_400_4);
  assign _zz_when_ArraySlice_l113_400_1 = (_zz_when_ArraySlice_l113_400_2 + _zz_when_ArraySlice_l113_400_3);
  assign _zz_when_ArraySlice_l113_400_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_400_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_400_4 = {1'd0, _zz_when_ArraySlice_l112_400};
  assign _zz__zz_when_ArraySlice_l173_400 = (_zz__zz_when_ArraySlice_l173_400_1 + _zz__zz_when_ArraySlice_l173_400_2);
  assign _zz__zz_when_ArraySlice_l173_400_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_400_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_400_3 = {1'd0, _zz_when_ArraySlice_l112_400};
  assign _zz_when_ArraySlice_l118_400_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_400 = _zz_when_ArraySlice_l118_400_1[5:0];
  assign _zz_when_ArraySlice_l173_400_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_400_2 = (_zz_when_ArraySlice_l173_400_3 + _zz_when_ArraySlice_l173_400_8);
  assign _zz_when_ArraySlice_l173_400_3 = (_zz_when_ArraySlice_l173_400 - _zz_when_ArraySlice_l173_400_4);
  assign _zz_when_ArraySlice_l173_400_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_400_6);
  assign _zz_when_ArraySlice_l173_400_4 = {1'd0, _zz_when_ArraySlice_l173_400_5};
  assign _zz_when_ArraySlice_l173_400_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_400_6 = {3'd0, _zz_when_ArraySlice_l173_400_7};
  assign _zz_when_ArraySlice_l173_400_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_401 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_401_1);
  assign _zz_when_ArraySlice_l165_401_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_401_1 = {2'd0, _zz_when_ArraySlice_l165_401_2};
  assign _zz_when_ArraySlice_l166_401 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_401_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_401_2);
  assign _zz_when_ArraySlice_l166_401_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_401_3);
  assign _zz_when_ArraySlice_l166_401_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_401_3 = {2'd0, _zz_when_ArraySlice_l166_401_4};
  assign _zz__zz_when_ArraySlice_l112_401 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_401 = (_zz_when_ArraySlice_l113_401_1 - _zz_when_ArraySlice_l113_401_4);
  assign _zz_when_ArraySlice_l113_401_1 = (_zz_when_ArraySlice_l113_401_2 + _zz_when_ArraySlice_l113_401_3);
  assign _zz_when_ArraySlice_l113_401_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_401_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_401_4 = {1'd0, _zz_when_ArraySlice_l112_401};
  assign _zz__zz_when_ArraySlice_l173_401 = (_zz__zz_when_ArraySlice_l173_401_1 + _zz__zz_when_ArraySlice_l173_401_2);
  assign _zz__zz_when_ArraySlice_l173_401_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_401_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_401_3 = {1'd0, _zz_when_ArraySlice_l112_401};
  assign _zz_when_ArraySlice_l118_401_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_401 = _zz_when_ArraySlice_l118_401_1[5:0];
  assign _zz_when_ArraySlice_l173_401_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_401_1 = {1'd0, _zz_when_ArraySlice_l173_401_2};
  assign _zz_when_ArraySlice_l173_401_3 = (_zz_when_ArraySlice_l173_401_4 + _zz_when_ArraySlice_l173_401_9);
  assign _zz_when_ArraySlice_l173_401_4 = (_zz_when_ArraySlice_l173_401 - _zz_when_ArraySlice_l173_401_5);
  assign _zz_when_ArraySlice_l173_401_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_401_7);
  assign _zz_when_ArraySlice_l173_401_5 = {1'd0, _zz_when_ArraySlice_l173_401_6};
  assign _zz_when_ArraySlice_l173_401_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_401_7 = {2'd0, _zz_when_ArraySlice_l173_401_8};
  assign _zz_when_ArraySlice_l173_401_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_402 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_402_1);
  assign _zz_when_ArraySlice_l165_402_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_402_1 = {1'd0, _zz_when_ArraySlice_l165_402_2};
  assign _zz_when_ArraySlice_l166_402 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_402_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_402_2);
  assign _zz_when_ArraySlice_l166_402_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_402_3);
  assign _zz_when_ArraySlice_l166_402_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_402_3 = {1'd0, _zz_when_ArraySlice_l166_402_4};
  assign _zz__zz_when_ArraySlice_l112_402 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_402 = (_zz_when_ArraySlice_l113_402_1 - _zz_when_ArraySlice_l113_402_4);
  assign _zz_when_ArraySlice_l113_402_1 = (_zz_when_ArraySlice_l113_402_2 + _zz_when_ArraySlice_l113_402_3);
  assign _zz_when_ArraySlice_l113_402_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_402_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_402_4 = {1'd0, _zz_when_ArraySlice_l112_402};
  assign _zz__zz_when_ArraySlice_l173_402 = (_zz__zz_when_ArraySlice_l173_402_1 + _zz__zz_when_ArraySlice_l173_402_2);
  assign _zz__zz_when_ArraySlice_l173_402_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_402_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_402_3 = {1'd0, _zz_when_ArraySlice_l112_402};
  assign _zz_when_ArraySlice_l118_402_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_402 = _zz_when_ArraySlice_l118_402_1[5:0];
  assign _zz_when_ArraySlice_l173_402_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_402_1 = {1'd0, _zz_when_ArraySlice_l173_402_2};
  assign _zz_when_ArraySlice_l173_402_3 = (_zz_when_ArraySlice_l173_402_4 + _zz_when_ArraySlice_l173_402_9);
  assign _zz_when_ArraySlice_l173_402_4 = (_zz_when_ArraySlice_l173_402 - _zz_when_ArraySlice_l173_402_5);
  assign _zz_when_ArraySlice_l173_402_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_402_7);
  assign _zz_when_ArraySlice_l173_402_5 = {1'd0, _zz_when_ArraySlice_l173_402_6};
  assign _zz_when_ArraySlice_l173_402_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_402_7 = {1'd0, _zz_when_ArraySlice_l173_402_8};
  assign _zz_when_ArraySlice_l173_402_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_403 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_403_1);
  assign _zz_when_ArraySlice_l165_403_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_403_1 = {1'd0, _zz_when_ArraySlice_l165_403_2};
  assign _zz_when_ArraySlice_l166_403 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_403_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_403_2);
  assign _zz_when_ArraySlice_l166_403_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_403_3);
  assign _zz_when_ArraySlice_l166_403_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_403_3 = {1'd0, _zz_when_ArraySlice_l166_403_4};
  assign _zz__zz_when_ArraySlice_l112_403 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_403 = (_zz_when_ArraySlice_l113_403_1 - _zz_when_ArraySlice_l113_403_4);
  assign _zz_when_ArraySlice_l113_403_1 = (_zz_when_ArraySlice_l113_403_2 + _zz_when_ArraySlice_l113_403_3);
  assign _zz_when_ArraySlice_l113_403_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_403_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_403_4 = {1'd0, _zz_when_ArraySlice_l112_403};
  assign _zz__zz_when_ArraySlice_l173_403 = (_zz__zz_when_ArraySlice_l173_403_1 + _zz__zz_when_ArraySlice_l173_403_2);
  assign _zz__zz_when_ArraySlice_l173_403_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_403_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_403_3 = {1'd0, _zz_when_ArraySlice_l112_403};
  assign _zz_when_ArraySlice_l118_403_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_403 = _zz_when_ArraySlice_l118_403_1[5:0];
  assign _zz_when_ArraySlice_l173_403_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_403_1 = {1'd0, _zz_when_ArraySlice_l173_403_2};
  assign _zz_when_ArraySlice_l173_403_3 = (_zz_when_ArraySlice_l173_403_4 + _zz_when_ArraySlice_l173_403_9);
  assign _zz_when_ArraySlice_l173_403_4 = (_zz_when_ArraySlice_l173_403 - _zz_when_ArraySlice_l173_403_5);
  assign _zz_when_ArraySlice_l173_403_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_403_7);
  assign _zz_when_ArraySlice_l173_403_5 = {1'd0, _zz_when_ArraySlice_l173_403_6};
  assign _zz_when_ArraySlice_l173_403_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_403_7 = {1'd0, _zz_when_ArraySlice_l173_403_8};
  assign _zz_when_ArraySlice_l173_403_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_404 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_404_1);
  assign _zz_when_ArraySlice_l165_404_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_404 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_404_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_404_2);
  assign _zz_when_ArraySlice_l166_404_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_404_3);
  assign _zz_when_ArraySlice_l166_404_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_404 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_404 = (_zz_when_ArraySlice_l113_404_1 - _zz_when_ArraySlice_l113_404_4);
  assign _zz_when_ArraySlice_l113_404_1 = (_zz_when_ArraySlice_l113_404_2 + _zz_when_ArraySlice_l113_404_3);
  assign _zz_when_ArraySlice_l113_404_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_404_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_404_4 = {1'd0, _zz_when_ArraySlice_l112_404};
  assign _zz__zz_when_ArraySlice_l173_404 = (_zz__zz_when_ArraySlice_l173_404_1 + _zz__zz_when_ArraySlice_l173_404_2);
  assign _zz__zz_when_ArraySlice_l173_404_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_404_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_404_3 = {1'd0, _zz_when_ArraySlice_l112_404};
  assign _zz_when_ArraySlice_l118_404_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_404 = _zz_when_ArraySlice_l118_404_1[5:0];
  assign _zz_when_ArraySlice_l173_404_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_404_1 = {1'd0, _zz_when_ArraySlice_l173_404_2};
  assign _zz_when_ArraySlice_l173_404_3 = (_zz_when_ArraySlice_l173_404_4 + _zz_when_ArraySlice_l173_404_8);
  assign _zz_when_ArraySlice_l173_404_4 = (_zz_when_ArraySlice_l173_404 - _zz_when_ArraySlice_l173_404_5);
  assign _zz_when_ArraySlice_l173_404_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_404_7);
  assign _zz_when_ArraySlice_l173_404_5 = {1'd0, _zz_when_ArraySlice_l173_404_6};
  assign _zz_when_ArraySlice_l173_404_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_404_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_405 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_405_1);
  assign _zz_when_ArraySlice_l165_405_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_405_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_405 = {1'd0, _zz_when_ArraySlice_l166_405_1};
  assign _zz_when_ArraySlice_l166_405_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_405_3);
  assign _zz_when_ArraySlice_l166_405_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_405_4);
  assign _zz_when_ArraySlice_l166_405_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_405 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_405 = (_zz_when_ArraySlice_l113_405_1 - _zz_when_ArraySlice_l113_405_4);
  assign _zz_when_ArraySlice_l113_405_1 = (_zz_when_ArraySlice_l113_405_2 + _zz_when_ArraySlice_l113_405_3);
  assign _zz_when_ArraySlice_l113_405_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_405_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_405_4 = {1'd0, _zz_when_ArraySlice_l112_405};
  assign _zz__zz_when_ArraySlice_l173_405 = (_zz__zz_when_ArraySlice_l173_405_1 + _zz__zz_when_ArraySlice_l173_405_2);
  assign _zz__zz_when_ArraySlice_l173_405_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_405_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_405_3 = {1'd0, _zz_when_ArraySlice_l112_405};
  assign _zz_when_ArraySlice_l118_405_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_405 = _zz_when_ArraySlice_l118_405_1[5:0];
  assign _zz_when_ArraySlice_l173_405_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_405_1 = {2'd0, _zz_when_ArraySlice_l173_405_2};
  assign _zz_when_ArraySlice_l173_405_3 = (_zz_when_ArraySlice_l173_405_4 + _zz_when_ArraySlice_l173_405_8);
  assign _zz_when_ArraySlice_l173_405_4 = (_zz_when_ArraySlice_l173_405 - _zz_when_ArraySlice_l173_405_5);
  assign _zz_when_ArraySlice_l173_405_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_405_7);
  assign _zz_when_ArraySlice_l173_405_5 = {1'd0, _zz_when_ArraySlice_l173_405_6};
  assign _zz_when_ArraySlice_l173_405_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_405_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_406 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_406_1);
  assign _zz_when_ArraySlice_l165_406_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_406_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_406 = {1'd0, _zz_when_ArraySlice_l166_406_1};
  assign _zz_when_ArraySlice_l166_406_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_406_3);
  assign _zz_when_ArraySlice_l166_406_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_406_4);
  assign _zz_when_ArraySlice_l166_406_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_406 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_406 = (_zz_when_ArraySlice_l113_406_1 - _zz_when_ArraySlice_l113_406_4);
  assign _zz_when_ArraySlice_l113_406_1 = (_zz_when_ArraySlice_l113_406_2 + _zz_when_ArraySlice_l113_406_3);
  assign _zz_when_ArraySlice_l113_406_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_406_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_406_4 = {1'd0, _zz_when_ArraySlice_l112_406};
  assign _zz__zz_when_ArraySlice_l173_406 = (_zz__zz_when_ArraySlice_l173_406_1 + _zz__zz_when_ArraySlice_l173_406_2);
  assign _zz__zz_when_ArraySlice_l173_406_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_406_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_406_3 = {1'd0, _zz_when_ArraySlice_l112_406};
  assign _zz_when_ArraySlice_l118_406_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_406 = _zz_when_ArraySlice_l118_406_1[5:0];
  assign _zz_when_ArraySlice_l173_406_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_406_1 = {2'd0, _zz_when_ArraySlice_l173_406_2};
  assign _zz_when_ArraySlice_l173_406_3 = (_zz_when_ArraySlice_l173_406_4 + _zz_when_ArraySlice_l173_406_8);
  assign _zz_when_ArraySlice_l173_406_4 = (_zz_when_ArraySlice_l173_406 - _zz_when_ArraySlice_l173_406_5);
  assign _zz_when_ArraySlice_l173_406_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_406_7);
  assign _zz_when_ArraySlice_l173_406_5 = {1'd0, _zz_when_ArraySlice_l173_406_6};
  assign _zz_when_ArraySlice_l173_406_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_406_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_407 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_407_1);
  assign _zz_when_ArraySlice_l165_407_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_407_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_407 = {2'd0, _zz_when_ArraySlice_l166_407_1};
  assign _zz_when_ArraySlice_l166_407_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_407_3);
  assign _zz_when_ArraySlice_l166_407_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_407_4);
  assign _zz_when_ArraySlice_l166_407_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_407 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_407 = (_zz_when_ArraySlice_l113_407_1 - _zz_when_ArraySlice_l113_407_4);
  assign _zz_when_ArraySlice_l113_407_1 = (_zz_when_ArraySlice_l113_407_2 + _zz_when_ArraySlice_l113_407_3);
  assign _zz_when_ArraySlice_l113_407_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_407_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_407_4 = {1'd0, _zz_when_ArraySlice_l112_407};
  assign _zz__zz_when_ArraySlice_l173_407 = (_zz__zz_when_ArraySlice_l173_407_1 + _zz__zz_when_ArraySlice_l173_407_2);
  assign _zz__zz_when_ArraySlice_l173_407_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_407_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_407_3 = {1'd0, _zz_when_ArraySlice_l112_407};
  assign _zz_when_ArraySlice_l118_407_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_407 = _zz_when_ArraySlice_l118_407_1[5:0];
  assign _zz_when_ArraySlice_l173_407_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_407_1 = {3'd0, _zz_when_ArraySlice_l173_407_2};
  assign _zz_when_ArraySlice_l173_407_3 = (_zz_when_ArraySlice_l173_407_4 + _zz_when_ArraySlice_l173_407_8);
  assign _zz_when_ArraySlice_l173_407_4 = (_zz_when_ArraySlice_l173_407 - _zz_when_ArraySlice_l173_407_5);
  assign _zz_when_ArraySlice_l173_407_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_407_7);
  assign _zz_when_ArraySlice_l173_407_5 = {1'd0, _zz_when_ArraySlice_l173_407_6};
  assign _zz_when_ArraySlice_l173_407_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_407_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_408 = (selectReadFifo_0 + _zz_when_ArraySlice_l165_408_1);
  assign _zz_when_ArraySlice_l165_408_2 = 3'b000;
  assign _zz_when_ArraySlice_l165_408_1 = {3'd0, _zz_when_ArraySlice_l165_408_2};
  assign _zz_when_ArraySlice_l166_408 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_408_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_408_3);
  assign _zz_when_ArraySlice_l166_408_1 = {1'd0, _zz_when_ArraySlice_l166_408_2};
  assign _zz_when_ArraySlice_l166_408_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_408_4);
  assign _zz_when_ArraySlice_l166_408_5 = 3'b000;
  assign _zz_when_ArraySlice_l166_408_4 = {3'd0, _zz_when_ArraySlice_l166_408_5};
  assign _zz__zz_when_ArraySlice_l112_408 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_408 = (_zz_when_ArraySlice_l113_408_1 - _zz_when_ArraySlice_l113_408_4);
  assign _zz_when_ArraySlice_l113_408_1 = (_zz_when_ArraySlice_l113_408_2 + _zz_when_ArraySlice_l113_408_3);
  assign _zz_when_ArraySlice_l113_408_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_408_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_408_4 = {1'd0, _zz_when_ArraySlice_l112_408};
  assign _zz__zz_when_ArraySlice_l173_408 = (_zz__zz_when_ArraySlice_l173_408_1 + _zz__zz_when_ArraySlice_l173_408_2);
  assign _zz__zz_when_ArraySlice_l173_408_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_408_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_408_3 = {1'd0, _zz_when_ArraySlice_l112_408};
  assign _zz_when_ArraySlice_l118_408_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_408 = _zz_when_ArraySlice_l118_408_1[5:0];
  assign _zz_when_ArraySlice_l173_408_1 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l173_408_2 = (_zz_when_ArraySlice_l173_408_3 + _zz_when_ArraySlice_l173_408_8);
  assign _zz_when_ArraySlice_l173_408_3 = (_zz_when_ArraySlice_l173_408 - _zz_when_ArraySlice_l173_408_4);
  assign _zz_when_ArraySlice_l173_408_5 = (selectReadFifo_0 + _zz_when_ArraySlice_l173_408_6);
  assign _zz_when_ArraySlice_l173_408_4 = {1'd0, _zz_when_ArraySlice_l173_408_5};
  assign _zz_when_ArraySlice_l173_408_7 = 3'b000;
  assign _zz_when_ArraySlice_l173_408_6 = {3'd0, _zz_when_ArraySlice_l173_408_7};
  assign _zz_when_ArraySlice_l173_408_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_409 = (selectReadFifo_1 + _zz_when_ArraySlice_l165_409_1);
  assign _zz_when_ArraySlice_l165_409_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l165_409_1 = {2'd0, _zz_when_ArraySlice_l165_409_2};
  assign _zz_when_ArraySlice_l166_409 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_409_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_409_2);
  assign _zz_when_ArraySlice_l166_409_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_409_3);
  assign _zz_when_ArraySlice_l166_409_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_409_3 = {2'd0, _zz_when_ArraySlice_l166_409_4};
  assign _zz__zz_when_ArraySlice_l112_409 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_409 = (_zz_when_ArraySlice_l113_409_1 - _zz_when_ArraySlice_l113_409_4);
  assign _zz_when_ArraySlice_l113_409_1 = (_zz_when_ArraySlice_l113_409_2 + _zz_when_ArraySlice_l113_409_3);
  assign _zz_when_ArraySlice_l113_409_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_409_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_409_4 = {1'd0, _zz_when_ArraySlice_l112_409};
  assign _zz__zz_when_ArraySlice_l173_409 = (_zz__zz_when_ArraySlice_l173_409_1 + _zz__zz_when_ArraySlice_l173_409_2);
  assign _zz__zz_when_ArraySlice_l173_409_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_409_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_409_3 = {1'd0, _zz_when_ArraySlice_l112_409};
  assign _zz_when_ArraySlice_l118_409_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_409 = _zz_when_ArraySlice_l118_409_1[5:0];
  assign _zz_when_ArraySlice_l173_409_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l173_409_1 = {1'd0, _zz_when_ArraySlice_l173_409_2};
  assign _zz_when_ArraySlice_l173_409_3 = (_zz_when_ArraySlice_l173_409_4 + _zz_when_ArraySlice_l173_409_9);
  assign _zz_when_ArraySlice_l173_409_4 = (_zz_when_ArraySlice_l173_409 - _zz_when_ArraySlice_l173_409_5);
  assign _zz_when_ArraySlice_l173_409_6 = (selectReadFifo_1 + _zz_when_ArraySlice_l173_409_7);
  assign _zz_when_ArraySlice_l173_409_5 = {1'd0, _zz_when_ArraySlice_l173_409_6};
  assign _zz_when_ArraySlice_l173_409_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l173_409_7 = {2'd0, _zz_when_ArraySlice_l173_409_8};
  assign _zz_when_ArraySlice_l173_409_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_410 = (selectReadFifo_2 + _zz_when_ArraySlice_l165_410_1);
  assign _zz_when_ArraySlice_l165_410_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l165_410_1 = {1'd0, _zz_when_ArraySlice_l165_410_2};
  assign _zz_when_ArraySlice_l166_410 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_410_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_410_2);
  assign _zz_when_ArraySlice_l166_410_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_410_3);
  assign _zz_when_ArraySlice_l166_410_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_410_3 = {1'd0, _zz_when_ArraySlice_l166_410_4};
  assign _zz__zz_when_ArraySlice_l112_410 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_410 = (_zz_when_ArraySlice_l113_410_1 - _zz_when_ArraySlice_l113_410_4);
  assign _zz_when_ArraySlice_l113_410_1 = (_zz_when_ArraySlice_l113_410_2 + _zz_when_ArraySlice_l113_410_3);
  assign _zz_when_ArraySlice_l113_410_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_410_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_410_4 = {1'd0, _zz_when_ArraySlice_l112_410};
  assign _zz__zz_when_ArraySlice_l173_410 = (_zz__zz_when_ArraySlice_l173_410_1 + _zz__zz_when_ArraySlice_l173_410_2);
  assign _zz__zz_when_ArraySlice_l173_410_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_410_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_410_3 = {1'd0, _zz_when_ArraySlice_l112_410};
  assign _zz_when_ArraySlice_l118_410_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_410 = _zz_when_ArraySlice_l118_410_1[5:0];
  assign _zz_when_ArraySlice_l173_410_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l173_410_1 = {1'd0, _zz_when_ArraySlice_l173_410_2};
  assign _zz_when_ArraySlice_l173_410_3 = (_zz_when_ArraySlice_l173_410_4 + _zz_when_ArraySlice_l173_410_9);
  assign _zz_when_ArraySlice_l173_410_4 = (_zz_when_ArraySlice_l173_410 - _zz_when_ArraySlice_l173_410_5);
  assign _zz_when_ArraySlice_l173_410_6 = (selectReadFifo_2 + _zz_when_ArraySlice_l173_410_7);
  assign _zz_when_ArraySlice_l173_410_5 = {1'd0, _zz_when_ArraySlice_l173_410_6};
  assign _zz_when_ArraySlice_l173_410_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l173_410_7 = {1'd0, _zz_when_ArraySlice_l173_410_8};
  assign _zz_when_ArraySlice_l173_410_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_411 = (selectReadFifo_3 + _zz_when_ArraySlice_l165_411_1);
  assign _zz_when_ArraySlice_l165_411_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l165_411_1 = {1'd0, _zz_when_ArraySlice_l165_411_2};
  assign _zz_when_ArraySlice_l166_411 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_411_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_411_2);
  assign _zz_when_ArraySlice_l166_411_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_411_3);
  assign _zz_when_ArraySlice_l166_411_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_411_3 = {1'd0, _zz_when_ArraySlice_l166_411_4};
  assign _zz__zz_when_ArraySlice_l112_411 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_411 = (_zz_when_ArraySlice_l113_411_1 - _zz_when_ArraySlice_l113_411_4);
  assign _zz_when_ArraySlice_l113_411_1 = (_zz_when_ArraySlice_l113_411_2 + _zz_when_ArraySlice_l113_411_3);
  assign _zz_when_ArraySlice_l113_411_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_411_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_411_4 = {1'd0, _zz_when_ArraySlice_l112_411};
  assign _zz__zz_when_ArraySlice_l173_411 = (_zz__zz_when_ArraySlice_l173_411_1 + _zz__zz_when_ArraySlice_l173_411_2);
  assign _zz__zz_when_ArraySlice_l173_411_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_411_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_411_3 = {1'd0, _zz_when_ArraySlice_l112_411};
  assign _zz_when_ArraySlice_l118_411_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_411 = _zz_when_ArraySlice_l118_411_1[5:0];
  assign _zz_when_ArraySlice_l173_411_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l173_411_1 = {1'd0, _zz_when_ArraySlice_l173_411_2};
  assign _zz_when_ArraySlice_l173_411_3 = (_zz_when_ArraySlice_l173_411_4 + _zz_when_ArraySlice_l173_411_9);
  assign _zz_when_ArraySlice_l173_411_4 = (_zz_when_ArraySlice_l173_411 - _zz_when_ArraySlice_l173_411_5);
  assign _zz_when_ArraySlice_l173_411_6 = (selectReadFifo_3 + _zz_when_ArraySlice_l173_411_7);
  assign _zz_when_ArraySlice_l173_411_5 = {1'd0, _zz_when_ArraySlice_l173_411_6};
  assign _zz_when_ArraySlice_l173_411_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l173_411_7 = {1'd0, _zz_when_ArraySlice_l173_411_8};
  assign _zz_when_ArraySlice_l173_411_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_412 = (selectReadFifo_4 + _zz_when_ArraySlice_l165_412_1);
  assign _zz_when_ArraySlice_l165_412_1 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_412 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_412_1 = (selectWriteFifo - _zz_when_ArraySlice_l166_412_2);
  assign _zz_when_ArraySlice_l166_412_2 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_412_3);
  assign _zz_when_ArraySlice_l166_412_3 = (bReg * 3'b100);
  assign _zz__zz_when_ArraySlice_l112_412 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_412 = (_zz_when_ArraySlice_l113_412_1 - _zz_when_ArraySlice_l113_412_4);
  assign _zz_when_ArraySlice_l113_412_1 = (_zz_when_ArraySlice_l113_412_2 + _zz_when_ArraySlice_l113_412_3);
  assign _zz_when_ArraySlice_l113_412_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_412_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_412_4 = {1'd0, _zz_when_ArraySlice_l112_412};
  assign _zz__zz_when_ArraySlice_l173_412 = (_zz__zz_when_ArraySlice_l173_412_1 + _zz__zz_when_ArraySlice_l173_412_2);
  assign _zz__zz_when_ArraySlice_l173_412_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_412_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_412_3 = {1'd0, _zz_when_ArraySlice_l112_412};
  assign _zz_when_ArraySlice_l118_412_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_412 = _zz_when_ArraySlice_l118_412_1[5:0];
  assign _zz_when_ArraySlice_l173_412_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l173_412_1 = {1'd0, _zz_when_ArraySlice_l173_412_2};
  assign _zz_when_ArraySlice_l173_412_3 = (_zz_when_ArraySlice_l173_412_4 + _zz_when_ArraySlice_l173_412_8);
  assign _zz_when_ArraySlice_l173_412_4 = (_zz_when_ArraySlice_l173_412 - _zz_when_ArraySlice_l173_412_5);
  assign _zz_when_ArraySlice_l173_412_6 = (selectReadFifo_4 + _zz_when_ArraySlice_l173_412_7);
  assign _zz_when_ArraySlice_l173_412_5 = {1'd0, _zz_when_ArraySlice_l173_412_6};
  assign _zz_when_ArraySlice_l173_412_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l173_412_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_413 = (selectReadFifo_5 + _zz_when_ArraySlice_l165_413_1);
  assign _zz_when_ArraySlice_l165_413_1 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_413_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_413 = {1'd0, _zz_when_ArraySlice_l166_413_1};
  assign _zz_when_ArraySlice_l166_413_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_413_3);
  assign _zz_when_ArraySlice_l166_413_3 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_413_4);
  assign _zz_when_ArraySlice_l166_413_4 = (bReg * 3'b101);
  assign _zz__zz_when_ArraySlice_l112_413 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_413 = (_zz_when_ArraySlice_l113_413_1 - _zz_when_ArraySlice_l113_413_4);
  assign _zz_when_ArraySlice_l113_413_1 = (_zz_when_ArraySlice_l113_413_2 + _zz_when_ArraySlice_l113_413_3);
  assign _zz_when_ArraySlice_l113_413_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_413_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_413_4 = {1'd0, _zz_when_ArraySlice_l112_413};
  assign _zz__zz_when_ArraySlice_l173_413 = (_zz__zz_when_ArraySlice_l173_413_1 + _zz__zz_when_ArraySlice_l173_413_2);
  assign _zz__zz_when_ArraySlice_l173_413_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_413_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_413_3 = {1'd0, _zz_when_ArraySlice_l112_413};
  assign _zz_when_ArraySlice_l118_413_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_413 = _zz_when_ArraySlice_l118_413_1[5:0];
  assign _zz_when_ArraySlice_l173_413_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l173_413_1 = {2'd0, _zz_when_ArraySlice_l173_413_2};
  assign _zz_when_ArraySlice_l173_413_3 = (_zz_when_ArraySlice_l173_413_4 + _zz_when_ArraySlice_l173_413_8);
  assign _zz_when_ArraySlice_l173_413_4 = (_zz_when_ArraySlice_l173_413 - _zz_when_ArraySlice_l173_413_5);
  assign _zz_when_ArraySlice_l173_413_6 = (selectReadFifo_5 + _zz_when_ArraySlice_l173_413_7);
  assign _zz_when_ArraySlice_l173_413_5 = {1'd0, _zz_when_ArraySlice_l173_413_6};
  assign _zz_when_ArraySlice_l173_413_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l173_413_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_414 = (selectReadFifo_6 + _zz_when_ArraySlice_l165_414_1);
  assign _zz_when_ArraySlice_l165_414_1 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_414_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_414 = {1'd0, _zz_when_ArraySlice_l166_414_1};
  assign _zz_when_ArraySlice_l166_414_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_414_3);
  assign _zz_when_ArraySlice_l166_414_3 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_414_4);
  assign _zz_when_ArraySlice_l166_414_4 = (bReg * 3'b110);
  assign _zz__zz_when_ArraySlice_l112_414 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_414 = (_zz_when_ArraySlice_l113_414_1 - _zz_when_ArraySlice_l113_414_4);
  assign _zz_when_ArraySlice_l113_414_1 = (_zz_when_ArraySlice_l113_414_2 + _zz_when_ArraySlice_l113_414_3);
  assign _zz_when_ArraySlice_l113_414_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_414_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_414_4 = {1'd0, _zz_when_ArraySlice_l112_414};
  assign _zz__zz_when_ArraySlice_l173_414 = (_zz__zz_when_ArraySlice_l173_414_1 + _zz__zz_when_ArraySlice_l173_414_2);
  assign _zz__zz_when_ArraySlice_l173_414_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_414_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_414_3 = {1'd0, _zz_when_ArraySlice_l112_414};
  assign _zz_when_ArraySlice_l118_414_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_414 = _zz_when_ArraySlice_l118_414_1[5:0];
  assign _zz_when_ArraySlice_l173_414_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l173_414_1 = {2'd0, _zz_when_ArraySlice_l173_414_2};
  assign _zz_when_ArraySlice_l173_414_3 = (_zz_when_ArraySlice_l173_414_4 + _zz_when_ArraySlice_l173_414_8);
  assign _zz_when_ArraySlice_l173_414_4 = (_zz_when_ArraySlice_l173_414 - _zz_when_ArraySlice_l173_414_5);
  assign _zz_when_ArraySlice_l173_414_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l173_414_7);
  assign _zz_when_ArraySlice_l173_414_5 = {1'd0, _zz_when_ArraySlice_l173_414_6};
  assign _zz_when_ArraySlice_l173_414_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l173_414_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l165_415 = (selectReadFifo_7 + _zz_when_ArraySlice_l165_415_1);
  assign _zz_when_ArraySlice_l165_415_1 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_415_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_415 = {2'd0, _zz_when_ArraySlice_l166_415_1};
  assign _zz_when_ArraySlice_l166_415_2 = (selectWriteFifo - _zz_when_ArraySlice_l166_415_3);
  assign _zz_when_ArraySlice_l166_415_3 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_415_4);
  assign _zz_when_ArraySlice_l166_415_4 = (bReg * 3'b111);
  assign _zz__zz_when_ArraySlice_l112_415 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_415 = (_zz_when_ArraySlice_l113_415_1 - _zz_when_ArraySlice_l113_415_4);
  assign _zz_when_ArraySlice_l113_415_1 = (_zz_when_ArraySlice_l113_415_2 + _zz_when_ArraySlice_l113_415_3);
  assign _zz_when_ArraySlice_l113_415_2 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l113_415_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l113_415_4 = {1'd0, _zz_when_ArraySlice_l112_415};
  assign _zz__zz_when_ArraySlice_l173_415 = (_zz__zz_when_ArraySlice_l173_415_1 + _zz__zz_when_ArraySlice_l173_415_2);
  assign _zz__zz_when_ArraySlice_l173_415_1 = {1'd0, wReg};
  assign _zz__zz_when_ArraySlice_l173_415_2 = (bReg * 4'b1000);
  assign _zz__zz_when_ArraySlice_l173_415_3 = {1'd0, _zz_when_ArraySlice_l112_415};
  assign _zz_when_ArraySlice_l118_415_1 = 7'h40;
  assign _zz_when_ArraySlice_l118_415 = _zz_when_ArraySlice_l118_415_1[5:0];
  assign _zz_when_ArraySlice_l173_415_2 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l173_415_1 = {3'd0, _zz_when_ArraySlice_l173_415_2};
  assign _zz_when_ArraySlice_l173_415_3 = (_zz_when_ArraySlice_l173_415_4 + _zz_when_ArraySlice_l173_415_8);
  assign _zz_when_ArraySlice_l173_415_4 = (_zz_when_ArraySlice_l173_415 - _zz_when_ArraySlice_l173_415_5);
  assign _zz_when_ArraySlice_l173_415_6 = (selectReadFifo_7 + _zz_when_ArraySlice_l173_415_7);
  assign _zz_when_ArraySlice_l173_415_5 = {1'd0, _zz_when_ArraySlice_l173_415_6};
  assign _zz_when_ArraySlice_l173_415_7 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l173_415_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l189_8 = (selectReadFifo_0 - _zz_when_ArraySlice_l189_8_1);
  assign _zz_when_ArraySlice_l189_8_1 = (selectReadFifo_0 % bReg);
  assign _zz_when_ArraySlice_l189_9 = (selectReadFifo_1 - _zz_when_ArraySlice_l189_9_1);
  assign _zz_when_ArraySlice_l189_9_1 = (selectReadFifo_1 % bReg);
  assign _zz_when_ArraySlice_l189_10 = (selectReadFifo_2 - _zz_when_ArraySlice_l189_10_1);
  assign _zz_when_ArraySlice_l189_10_1 = (selectReadFifo_2 % bReg);
  assign _zz_when_ArraySlice_l189_11 = (selectReadFifo_3 - _zz_when_ArraySlice_l189_11_1);
  assign _zz_when_ArraySlice_l189_11_1 = (selectReadFifo_3 % bReg);
  assign _zz_when_ArraySlice_l189_12 = (selectReadFifo_4 - _zz_when_ArraySlice_l189_12_1);
  assign _zz_when_ArraySlice_l189_12_1 = (selectReadFifo_4 % bReg);
  assign _zz_when_ArraySlice_l189_13 = (selectReadFifo_5 - _zz_when_ArraySlice_l189_13_1);
  assign _zz_when_ArraySlice_l189_13_1 = (selectReadFifo_5 % bReg);
  assign _zz_when_ArraySlice_l189_14 = (selectReadFifo_6 - _zz_when_ArraySlice_l189_14_1);
  assign _zz_when_ArraySlice_l189_14_1 = (selectReadFifo_6 % bReg);
  assign _zz_when_ArraySlice_l189_15 = (selectReadFifo_7 - _zz_when_ArraySlice_l189_15_1);
  assign _zz_when_ArraySlice_l189_15_1 = (selectReadFifo_7 % bReg);
  assign _zz_when_ArraySlice_l189_16 = (selectReadFifo_0 - _zz_when_ArraySlice_l189_16_1);
  assign _zz_when_ArraySlice_l189_16_1 = (selectReadFifo_0 % bReg);
  assign _zz_when_ArraySlice_l189_17 = (selectReadFifo_1 - _zz_when_ArraySlice_l189_17_1);
  assign _zz_when_ArraySlice_l189_17_1 = (selectReadFifo_1 % bReg);
  assign _zz_when_ArraySlice_l189_18 = (selectReadFifo_2 - _zz_when_ArraySlice_l189_18_1);
  assign _zz_when_ArraySlice_l189_18_1 = (selectReadFifo_2 % bReg);
  assign _zz_when_ArraySlice_l189_19 = (selectReadFifo_3 - _zz_when_ArraySlice_l189_19_1);
  assign _zz_when_ArraySlice_l189_19_1 = (selectReadFifo_3 % bReg);
  assign _zz_when_ArraySlice_l189_20 = (selectReadFifo_4 - _zz_when_ArraySlice_l189_20_1);
  assign _zz_when_ArraySlice_l189_20_1 = (selectReadFifo_4 % bReg);
  assign _zz_when_ArraySlice_l189_21 = (selectReadFifo_5 - _zz_when_ArraySlice_l189_21_1);
  assign _zz_when_ArraySlice_l189_21_1 = (selectReadFifo_5 % bReg);
  assign _zz_when_ArraySlice_l189_22 = (selectReadFifo_6 - _zz_when_ArraySlice_l189_22_1);
  assign _zz_when_ArraySlice_l189_22_1 = (selectReadFifo_6 % bReg);
  assign _zz_when_ArraySlice_l189_23 = (selectReadFifo_7 - _zz_when_ArraySlice_l189_23_1);
  assign _zz_when_ArraySlice_l189_23_1 = (selectReadFifo_7 % bReg);
  assign _zz_when_ArraySlice_l398 = ((((holdReadOp_0 == _zz_when_ArraySlice_l398_1) && (holdReadOp_1 == _zz_when_ArraySlice_l398_2)) && (holdReadOp_2 == 1'b1)) && (holdReadOp_3 == 1'b1));
  assign _zz_when_ArraySlice_l398_3 = (holdReadOp_4 == 1'b1);
  assign _zz_when_ArraySlice_l398_4 = 1'b1;
  assign _zz_when_ArraySlice_l398_5 = ((((debug_0_1 == _zz_when_ArraySlice_l398_6) && (debug_1_1 == _zz_when_ArraySlice_l398_7)) && (debug_2_1 == 1'b1)) && (debug_3_1 == 1'b1));
  assign _zz_when_ArraySlice_l398_8 = (debug_4_1 == 1'b1);
  assign _zz_when_ArraySlice_l398_9 = 1'b1;
  assign _zz_when_ArraySlice_l398_1 = 1'b1;
  assign _zz_when_ArraySlice_l398_2 = 1'b1;
  assign _zz_when_ArraySlice_l398_6 = 1'b1;
  assign _zz_when_ArraySlice_l398_7 = 1'b1;
  assign _zz_when_ArraySlice_l418 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l418_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l418_2 = 1'b1;
  assign _zz_when_ArraySlice_l418_3 = (((debug_0_2 == 1'b1) && (debug_1_2 == 1'b1)) && (debug_2_2 == 1'b1));
  assign _zz_when_ArraySlice_l418_4 = (debug_3_2 == 1'b1);
  assign _zz_when_ArraySlice_l418_5 = 1'b1;
  assign _zz_when_ArraySlice_l444 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l444_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l444_2 = 1'b1;
  assign _zz_when_ArraySlice_l444_3 = (((debug_0_3 == 1'b1) && (debug_1_3 == 1'b1)) && (debug_2_3 == 1'b1));
  assign _zz_when_ArraySlice_l444_4 = (debug_3_3 == 1'b1);
  assign _zz_when_ArraySlice_l444_5 = 1'b1;
  assign _zz_when_ArraySlice_l398_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l398_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l398_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l398_1_4 = (((debug_0_4 == 1'b1) && (debug_1_4 == 1'b1)) && (debug_2_4 == 1'b1));
  assign _zz_when_ArraySlice_l398_1_5 = (debug_3_4 == 1'b1);
  assign _zz_when_ArraySlice_l398_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l418_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l418_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l418_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l418_1_4 = (((debug_0_5 == 1'b1) && (debug_1_5 == 1'b1)) && (debug_2_5 == 1'b1));
  assign _zz_when_ArraySlice_l418_1_5 = (debug_3_5 == 1'b1);
  assign _zz_when_ArraySlice_l418_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l444_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l444_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l444_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l444_1_4 = (((debug_0_6 == 1'b1) && (debug_1_6 == 1'b1)) && (debug_2_6 == 1'b1));
  assign _zz_when_ArraySlice_l444_1_5 = (debug_3_6 == 1'b1);
  assign _zz_when_ArraySlice_l444_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l398_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l398_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l398_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l398_2_4 = (((debug_0_7 == 1'b1) && (debug_1_7 == 1'b1)) && (debug_2_7 == 1'b1));
  assign _zz_when_ArraySlice_l398_2_5 = (debug_3_7 == 1'b1);
  assign _zz_when_ArraySlice_l398_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l418_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l418_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l418_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l418_2_4 = (((debug_0_8 == 1'b1) && (debug_1_8 == 1'b1)) && (debug_2_8 == 1'b1));
  assign _zz_when_ArraySlice_l418_2_5 = (debug_3_8 == 1'b1);
  assign _zz_when_ArraySlice_l418_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l444_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l444_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l444_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l444_2_4 = (((debug_0_9 == 1'b1) && (debug_1_9 == 1'b1)) && (debug_2_9 == 1'b1));
  assign _zz_when_ArraySlice_l444_2_5 = (debug_3_9 == 1'b1);
  assign _zz_when_ArraySlice_l444_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l398_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l398_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l398_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l398_3_4 = (((debug_0_10 == 1'b1) && (debug_1_10 == 1'b1)) && (debug_2_10 == 1'b1));
  assign _zz_when_ArraySlice_l398_3_5 = (debug_3_10 == 1'b1);
  assign _zz_when_ArraySlice_l398_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l418_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l418_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l418_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l418_3_4 = (((debug_0_11 == 1'b1) && (debug_1_11 == 1'b1)) && (debug_2_11 == 1'b1));
  assign _zz_when_ArraySlice_l418_3_5 = (debug_3_11 == 1'b1);
  assign _zz_when_ArraySlice_l418_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l444_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l444_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l444_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l444_3_4 = (((debug_0_12 == 1'b1) && (debug_1_12 == 1'b1)) && (debug_2_12 == 1'b1));
  assign _zz_when_ArraySlice_l444_3_5 = (debug_3_12 == 1'b1);
  assign _zz_when_ArraySlice_l444_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l398_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l398_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l398_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l398_4_4 = (((debug_0_13 == 1'b1) && (debug_1_13 == 1'b1)) && (debug_2_13 == 1'b1));
  assign _zz_when_ArraySlice_l398_4_5 = (debug_3_13 == 1'b1);
  assign _zz_when_ArraySlice_l398_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l418_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l418_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l418_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l418_4_4 = (((debug_0_14 == 1'b1) && (debug_1_14 == 1'b1)) && (debug_2_14 == 1'b1));
  assign _zz_when_ArraySlice_l418_4_5 = (debug_3_14 == 1'b1);
  assign _zz_when_ArraySlice_l418_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l444_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l444_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l444_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l444_4_4 = (((debug_0_15 == 1'b1) && (debug_1_15 == 1'b1)) && (debug_2_15 == 1'b1));
  assign _zz_when_ArraySlice_l444_4_5 = (debug_3_15 == 1'b1);
  assign _zz_when_ArraySlice_l444_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l398_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l398_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l398_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l398_5_4 = (((debug_0_16 == 1'b1) && (debug_1_16 == 1'b1)) && (debug_2_16 == 1'b1));
  assign _zz_when_ArraySlice_l398_5_5 = (debug_3_16 == 1'b1);
  assign _zz_when_ArraySlice_l398_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l418_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l418_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l418_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l418_5_4 = (((debug_0_17 == 1'b1) && (debug_1_17 == 1'b1)) && (debug_2_17 == 1'b1));
  assign _zz_when_ArraySlice_l418_5_5 = (debug_3_17 == 1'b1);
  assign _zz_when_ArraySlice_l418_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l444_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l444_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l444_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l444_5_4 = (((debug_0_18 == 1'b1) && (debug_1_18 == 1'b1)) && (debug_2_18 == 1'b1));
  assign _zz_when_ArraySlice_l444_5_5 = (debug_3_18 == 1'b1);
  assign _zz_when_ArraySlice_l444_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l398_6_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l398_6_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l398_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l398_6_4 = (((debug_0_19 == 1'b1) && (debug_1_19 == 1'b1)) && (debug_2_19 == 1'b1));
  assign _zz_when_ArraySlice_l398_6_5 = (debug_3_19 == 1'b1);
  assign _zz_when_ArraySlice_l398_6_6 = 1'b1;
  assign _zz_when_ArraySlice_l418_6 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l418_6_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l418_6_2 = 1'b1;
  assign _zz_when_ArraySlice_l418_6_3 = (((debug_0_20 == 1'b1) && (debug_1_20 == 1'b1)) && (debug_2_20 == 1'b1));
  assign _zz_when_ArraySlice_l418_6_4 = (debug_3_20 == 1'b1);
  assign _zz_when_ArraySlice_l418_6_5 = 1'b1;
  assign _zz_when_ArraySlice_l444_6 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l444_6_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l444_6_2 = 1'b1;
  assign _zz_when_ArraySlice_l444_6_3 = (((debug_0_21 == 1'b1) && (debug_1_21 == 1'b1)) && (debug_2_21 == 1'b1));
  assign _zz_when_ArraySlice_l444_6_4 = (debug_3_21 == 1'b1);
  assign _zz_when_ArraySlice_l444_6_5 = 1'b1;
  assign _zz_when_ArraySlice_l398_7_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l398_7_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l398_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l398_7_4 = (((debug_0_22 == 1'b1) && (debug_1_22 == 1'b1)) && (debug_2_22 == 1'b1));
  assign _zz_when_ArraySlice_l398_7_5 = (debug_3_22 == 1'b1);
  assign _zz_when_ArraySlice_l398_7_6 = 1'b1;
  assign _zz_when_ArraySlice_l418_7 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l418_7_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l418_7_2 = 1'b1;
  assign _zz_when_ArraySlice_l418_7_3 = (((debug_0_23 == 1'b1) && (debug_1_23 == 1'b1)) && (debug_2_23 == 1'b1));
  assign _zz_when_ArraySlice_l418_7_4 = (debug_3_23 == 1'b1);
  assign _zz_when_ArraySlice_l418_7_5 = 1'b1;
  assign _zz_when_ArraySlice_l444_7 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l444_7_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l444_7_2 = 1'b1;
  assign _zz_when_ArraySlice_l444_7_3 = (((debug_0_24 == 1'b1) && (debug_1_24 == 1'b1)) && (debug_2_24 == 1'b1));
  assign _zz_when_ArraySlice_l444_7_4 = (debug_3_24 == 1'b1);
  assign _zz_when_ArraySlice_l444_7_5 = 1'b1;
  assign _zz_when_ArraySlice_l465 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l465_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l465_2 = 1'b1;
  assign _zz_when_ArraySlice_l465_3 = (((debug_0_25 == 1'b1) && (debug_1_25 == 1'b1)) && (debug_2_25 == 1'b1));
  assign _zz_when_ArraySlice_l465_4 = (debug_3_25 == 1'b1);
  assign _zz_when_ArraySlice_l465_5 = 1'b1;
  assign _zz_when_ArraySlice_l265 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l265_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l265_2 = 1'b1;
  assign _zz_when_ArraySlice_l265_3 = (((debug_0_26 == 1'b1) && (debug_1_26 == 1'b1)) && (debug_2_26 == 1'b1));
  assign _zz_when_ArraySlice_l265_4 = (debug_3_26 == 1'b1);
  assign _zz_when_ArraySlice_l265_5 = 1'b1;
  assign _zz_when_ArraySlice_l285 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l285_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l285_2 = 1'b1;
  assign _zz_when_ArraySlice_l285_3 = (((debug_0_27 == 1'b1) && (debug_1_27 == 1'b1)) && (debug_2_27 == 1'b1));
  assign _zz_when_ArraySlice_l285_4 = (debug_3_27 == 1'b1);
  assign _zz_when_ArraySlice_l285_5 = 1'b1;
  assign _zz_when_ArraySlice_l311 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l311_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l311_2 = 1'b1;
  assign _zz_when_ArraySlice_l311_3 = (((debug_0_28 == 1'b1) && (debug_1_28 == 1'b1)) && (debug_2_28 == 1'b1));
  assign _zz_when_ArraySlice_l311_4 = (debug_3_28 == 1'b1);
  assign _zz_when_ArraySlice_l311_5 = 1'b1;
  assign _zz_when_ArraySlice_l265_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l265_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l265_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l265_1_4 = (((debug_0_29 == 1'b1) && (debug_1_29 == 1'b1)) && (debug_2_29 == 1'b1));
  assign _zz_when_ArraySlice_l265_1_5 = (debug_3_29 == 1'b1);
  assign _zz_when_ArraySlice_l265_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l285_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l285_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l285_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l285_1_4 = (((debug_0_30 == 1'b1) && (debug_1_30 == 1'b1)) && (debug_2_30 == 1'b1));
  assign _zz_when_ArraySlice_l285_1_5 = (debug_3_30 == 1'b1);
  assign _zz_when_ArraySlice_l285_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l311_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l311_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l311_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l311_1_4 = (((debug_0_31 == 1'b1) && (debug_1_31 == 1'b1)) && (debug_2_31 == 1'b1));
  assign _zz_when_ArraySlice_l311_1_5 = (debug_3_31 == 1'b1);
  assign _zz_when_ArraySlice_l311_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l265_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l265_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l265_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l265_2_4 = (((debug_0_32 == 1'b1) && (debug_1_32 == 1'b1)) && (debug_2_32 == 1'b1));
  assign _zz_when_ArraySlice_l265_2_5 = (debug_3_32 == 1'b1);
  assign _zz_when_ArraySlice_l265_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l285_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l285_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l285_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l285_2_4 = (((debug_0_33 == 1'b1) && (debug_1_33 == 1'b1)) && (debug_2_33 == 1'b1));
  assign _zz_when_ArraySlice_l285_2_5 = (debug_3_33 == 1'b1);
  assign _zz_when_ArraySlice_l285_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l311_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l311_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l311_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l311_2_4 = (((debug_0_34 == 1'b1) && (debug_1_34 == 1'b1)) && (debug_2_34 == 1'b1));
  assign _zz_when_ArraySlice_l311_2_5 = (debug_3_34 == 1'b1);
  assign _zz_when_ArraySlice_l311_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l265_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l265_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l265_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l265_3_4 = (((debug_0_35 == 1'b1) && (debug_1_35 == 1'b1)) && (debug_2_35 == 1'b1));
  assign _zz_when_ArraySlice_l265_3_5 = (debug_3_35 == 1'b1);
  assign _zz_when_ArraySlice_l265_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l285_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l285_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l285_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l285_3_4 = (((debug_0_36 == 1'b1) && (debug_1_36 == 1'b1)) && (debug_2_36 == 1'b1));
  assign _zz_when_ArraySlice_l285_3_5 = (debug_3_36 == 1'b1);
  assign _zz_when_ArraySlice_l285_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l311_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l311_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l311_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l311_3_4 = (((debug_0_37 == 1'b1) && (debug_1_37 == 1'b1)) && (debug_2_37 == 1'b1));
  assign _zz_when_ArraySlice_l311_3_5 = (debug_3_37 == 1'b1);
  assign _zz_when_ArraySlice_l311_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l265_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l265_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l265_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l265_4_4 = (((debug_0_38 == 1'b1) && (debug_1_38 == 1'b1)) && (debug_2_38 == 1'b1));
  assign _zz_when_ArraySlice_l265_4_5 = (debug_3_38 == 1'b1);
  assign _zz_when_ArraySlice_l265_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l285_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l285_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l285_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l285_4_4 = (((debug_0_39 == 1'b1) && (debug_1_39 == 1'b1)) && (debug_2_39 == 1'b1));
  assign _zz_when_ArraySlice_l285_4_5 = (debug_3_39 == 1'b1);
  assign _zz_when_ArraySlice_l285_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l311_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l311_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l311_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l311_4_4 = (((debug_0_40 == 1'b1) && (debug_1_40 == 1'b1)) && (debug_2_40 == 1'b1));
  assign _zz_when_ArraySlice_l311_4_5 = (debug_3_40 == 1'b1);
  assign _zz_when_ArraySlice_l311_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l265_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l265_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l265_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l265_5_4 = (((debug_0_41 == 1'b1) && (debug_1_41 == 1'b1)) && (debug_2_41 == 1'b1));
  assign _zz_when_ArraySlice_l265_5_5 = (debug_3_41 == 1'b1);
  assign _zz_when_ArraySlice_l265_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l285_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l285_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l285_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l285_5_4 = (((debug_0_42 == 1'b1) && (debug_1_42 == 1'b1)) && (debug_2_42 == 1'b1));
  assign _zz_when_ArraySlice_l285_5_5 = (debug_3_42 == 1'b1);
  assign _zz_when_ArraySlice_l285_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l311_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l311_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l311_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l311_5_4 = (((debug_0_43 == 1'b1) && (debug_1_43 == 1'b1)) && (debug_2_43 == 1'b1));
  assign _zz_when_ArraySlice_l311_5_5 = (debug_3_43 == 1'b1);
  assign _zz_when_ArraySlice_l311_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l265_6 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l265_6_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l265_6_2 = 1'b1;
  assign _zz_when_ArraySlice_l265_6_3 = (((debug_0_44 == 1'b1) && (debug_1_44 == 1'b1)) && (debug_2_44 == 1'b1));
  assign _zz_when_ArraySlice_l265_6_4 = (debug_3_44 == 1'b1);
  assign _zz_when_ArraySlice_l265_6_5 = 1'b1;
  assign _zz_when_ArraySlice_l285_6 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l285_6_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l285_6_2 = 1'b1;
  assign _zz_when_ArraySlice_l285_6_3 = (((debug_0_45 == 1'b1) && (debug_1_45 == 1'b1)) && (debug_2_45 == 1'b1));
  assign _zz_when_ArraySlice_l285_6_4 = (debug_3_45 == 1'b1);
  assign _zz_when_ArraySlice_l285_6_5 = 1'b1;
  assign _zz_when_ArraySlice_l311_6 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l311_6_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l311_6_2 = 1'b1;
  assign _zz_when_ArraySlice_l311_6_3 = (((debug_0_46 == 1'b1) && (debug_1_46 == 1'b1)) && (debug_2_46 == 1'b1));
  assign _zz_when_ArraySlice_l311_6_4 = (debug_3_46 == 1'b1);
  assign _zz_when_ArraySlice_l311_6_5 = 1'b1;
  assign _zz_when_ArraySlice_l265_7 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l265_7_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l265_7_2 = 1'b1;
  assign _zz_when_ArraySlice_l265_7_3 = (((debug_0_47 == 1'b1) && (debug_1_47 == 1'b1)) && (debug_2_47 == 1'b1));
  assign _zz_when_ArraySlice_l265_7_4 = (debug_3_47 == 1'b1);
  assign _zz_when_ArraySlice_l265_7_5 = 1'b1;
  assign _zz_when_ArraySlice_l285_7 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l285_7_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l285_7_2 = 1'b1;
  assign _zz_when_ArraySlice_l285_7_3 = (((debug_0_48 == 1'b1) && (debug_1_48 == 1'b1)) && (debug_2_48 == 1'b1));
  assign _zz_when_ArraySlice_l285_7_4 = (debug_3_48 == 1'b1);
  assign _zz_when_ArraySlice_l285_7_5 = 1'b1;
  assign _zz_when_ArraySlice_l311_7 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l311_7_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l311_7_2 = 1'b1;
  assign _zz_when_ArraySlice_l311_7_3 = (((debug_0_49 == 1'b1) && (debug_1_49 == 1'b1)) && (debug_2_49 == 1'b1));
  assign _zz_when_ArraySlice_l311_7_4 = (debug_3_49 == 1'b1);
  assign _zz_when_ArraySlice_l311_7_5 = 1'b1;
  assign _zz_when_ArraySlice_l333_8 = 1'b0;
  assign _zz_when_ArraySlice_l333_9 = 1'b0;
  assign _zz_when_ArraySlice_l350 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l350_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l350_2 = 1'b1;
  assign _zz_when_ArraySlice_l350_3 = (((debug_0_50 == 1'b1) && (debug_1_50 == 1'b1)) && (debug_2_50 == 1'b1));
  assign _zz_when_ArraySlice_l350_4 = (debug_3_50 == 1'b1);
  assign _zz_when_ArraySlice_l350_5 = 1'b1;
  assign _zz_when_ArraySlice_l354_8 = (((_zz_when_ArraySlice_l354_9 && _zz_when_ArraySlice_l354_10) && (holdReadOp_3 == _zz_when_ArraySlice_l354_11)) && (holdReadOp_4 == 1'b1));
  assign _zz_when_ArraySlice_l354_12 = (holdReadOp_5 == 1'b1);
  assign _zz_when_ArraySlice_l354_13 = 1'b1;
  assign _zz_when_ArraySlice_l354_14 = (((_zz_when_ArraySlice_l354_15 && _zz_when_ArraySlice_l354_16) && (debug_4_51 == _zz_when_ArraySlice_l354_17)) && (debug_5_51 == 1'b1));
  assign _zz_when_ArraySlice_l354_18 = (debug_6_51 == 1'b1);
  assign _zz_when_ArraySlice_l354_19 = 1'b1;
  assign _zz_when_ArraySlice_l354_20 = (((_zz_when_ArraySlice_l354_21 || _zz_when_ArraySlice_l354_22) || (_zz_when_ArraySlice_l354_3 != _zz_when_ArraySlice_l354_23)) || (_zz_when_ArraySlice_l354_4 != 1'b0));
  assign _zz_when_ArraySlice_l354_24 = (_zz_when_ArraySlice_l354_5 != 1'b0);
  assign _zz_when_ArraySlice_l354_25 = 1'b0;
  assign _zz_when_ArraySlice_l354_9 = ((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1));
  assign _zz_when_ArraySlice_l354_10 = (holdReadOp_2 == 1'b1);
  assign _zz_when_ArraySlice_l354_11 = 1'b1;
  assign _zz_when_ArraySlice_l354_15 = (((debug_0_51 == 1'b1) && (debug_1_51 == 1'b1)) && (debug_2_51 == 1'b1));
  assign _zz_when_ArraySlice_l354_16 = (debug_3_51 == 1'b1);
  assign _zz_when_ArraySlice_l354_17 = 1'b1;
  assign _zz_when_ArraySlice_l354_21 = ((_zz_when_ArraySlice_l354 != 1'b0) || (_zz_when_ArraySlice_l354_1 != 1'b0));
  assign _zz_when_ArraySlice_l354_22 = (_zz_when_ArraySlice_l354_2 != 1'b0);
  assign _zz_when_ArraySlice_l354_23 = 1'b0;
  StreamFifo fifoGroup_0 (
    .io_push_valid      (fifoGroup_0_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_0_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_0_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_0_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_0_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_0_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                               ), //i
    .io_occupancy       (fifoGroup_0_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_0_io_availability[6:0]   ), //o
    .clk                (clk                                ), //i
    .resetn             (resetn                             )  //i
  );
  StreamFifo fifoGroup_1 (
    .io_push_valid      (fifoGroup_1_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_1_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_1_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_1_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_1_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_1_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                               ), //i
    .io_occupancy       (fifoGroup_1_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_1_io_availability[6:0]   ), //o
    .clk                (clk                                ), //i
    .resetn             (resetn                             )  //i
  );
  StreamFifo fifoGroup_2 (
    .io_push_valid      (fifoGroup_2_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_2_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_2_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_2_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_2_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_2_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                               ), //i
    .io_occupancy       (fifoGroup_2_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_2_io_availability[6:0]   ), //o
    .clk                (clk                                ), //i
    .resetn             (resetn                             )  //i
  );
  StreamFifo fifoGroup_3 (
    .io_push_valid      (fifoGroup_3_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_3_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_3_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_3_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_3_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_3_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                               ), //i
    .io_occupancy       (fifoGroup_3_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_3_io_availability[6:0]   ), //o
    .clk                (clk                                ), //i
    .resetn             (resetn                             )  //i
  );
  StreamFifo fifoGroup_4 (
    .io_push_valid      (fifoGroup_4_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_4_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_4_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_4_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_4_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_4_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                               ), //i
    .io_occupancy       (fifoGroup_4_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_4_io_availability[6:0]   ), //o
    .clk                (clk                                ), //i
    .resetn             (resetn                             )  //i
  );
  StreamFifo fifoGroup_5 (
    .io_push_valid      (fifoGroup_5_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_5_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_5_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_5_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_5_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_5_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                               ), //i
    .io_occupancy       (fifoGroup_5_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_5_io_availability[6:0]   ), //o
    .clk                (clk                                ), //i
    .resetn             (resetn                             )  //i
  );
  StreamFifo fifoGroup_6 (
    .io_push_valid      (fifoGroup_6_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_6_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_6_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_6_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_6_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_6_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                               ), //i
    .io_occupancy       (fifoGroup_6_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_6_io_availability[6:0]   ), //o
    .clk                (clk                                ), //i
    .resetn             (resetn                             )  //i
  );
  StreamFifo fifoGroup_7 (
    .io_push_valid      (fifoGroup_7_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_7_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_7_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_7_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_7_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_7_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                               ), //i
    .io_occupancy       (fifoGroup_7_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_7_io_availability[6:0]   ), //o
    .clk                (clk                                ), //i
    .resetn             (resetn                             )  //i
  );
  StreamFifo fifoGroup_8 (
    .io_push_valid      (fifoGroup_8_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_8_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_8_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_8_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_8_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_8_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                               ), //i
    .io_occupancy       (fifoGroup_8_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_8_io_availability[6:0]   ), //o
    .clk                (clk                                ), //i
    .resetn             (resetn                             )  //i
  );
  StreamFifo fifoGroup_9 (
    .io_push_valid      (fifoGroup_9_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_9_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_9_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_9_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_9_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_9_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                               ), //i
    .io_occupancy       (fifoGroup_9_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_9_io_availability[6:0]   ), //o
    .clk                (clk                                ), //i
    .resetn             (resetn                             )  //i
  );
  StreamFifo fifoGroup_10 (
    .io_push_valid      (fifoGroup_10_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_10_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_10_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_10_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_10_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_10_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_10_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_10_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_11 (
    .io_push_valid      (fifoGroup_11_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_11_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_11_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_11_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_11_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_11_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_11_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_11_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_12 (
    .io_push_valid      (fifoGroup_12_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_12_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_12_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_12_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_12_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_12_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_12_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_12_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_13 (
    .io_push_valid      (fifoGroup_13_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_13_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_13_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_13_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_13_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_13_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_13_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_13_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_14 (
    .io_push_valid      (fifoGroup_14_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_14_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_14_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_14_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_14_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_14_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_14_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_14_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_15 (
    .io_push_valid      (fifoGroup_15_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_15_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_15_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_15_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_15_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_15_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_15_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_15_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_16 (
    .io_push_valid      (fifoGroup_16_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_16_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_16_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_16_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_16_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_16_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_16_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_16_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_17 (
    .io_push_valid      (fifoGroup_17_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_17_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_17_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_17_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_17_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_17_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_17_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_17_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_18 (
    .io_push_valid      (fifoGroup_18_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_18_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_18_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_18_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_18_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_18_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_18_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_18_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_19 (
    .io_push_valid      (fifoGroup_19_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_19_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_19_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_19_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_19_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_19_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_19_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_19_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_20 (
    .io_push_valid      (fifoGroup_20_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_20_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_20_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_20_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_20_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_20_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_20_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_20_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_21 (
    .io_push_valid      (fifoGroup_21_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_21_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_21_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_21_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_21_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_21_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_21_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_21_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_22 (
    .io_push_valid      (fifoGroup_22_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_22_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_22_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_22_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_22_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_22_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_22_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_22_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_23 (
    .io_push_valid      (fifoGroup_23_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_23_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_23_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_23_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_23_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_23_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_23_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_23_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_24 (
    .io_push_valid      (fifoGroup_24_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_24_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_24_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_24_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_24_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_24_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_24_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_24_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_25 (
    .io_push_valid      (fifoGroup_25_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_25_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_25_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_25_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_25_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_25_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_25_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_25_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_26 (
    .io_push_valid      (fifoGroup_26_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_26_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_26_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_26_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_26_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_26_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_26_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_26_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_27 (
    .io_push_valid      (fifoGroup_27_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_27_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_27_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_27_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_27_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_27_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_27_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_27_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_28 (
    .io_push_valid      (fifoGroup_28_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_28_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_28_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_28_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_28_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_28_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_28_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_28_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_29 (
    .io_push_valid      (fifoGroup_29_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_29_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_29_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_29_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_29_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_29_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_29_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_29_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_30 (
    .io_push_valid      (fifoGroup_30_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_30_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_30_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_30_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_30_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_30_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_30_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_30_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_31 (
    .io_push_valid      (fifoGroup_31_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_31_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_31_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_31_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_31_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_31_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_31_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_31_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_32 (
    .io_push_valid      (fifoGroup_32_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_32_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_32_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_32_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_32_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_32_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_32_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_32_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_33 (
    .io_push_valid      (fifoGroup_33_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_33_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_33_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_33_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_33_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_33_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_33_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_33_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_34 (
    .io_push_valid      (fifoGroup_34_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_34_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_34_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_34_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_34_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_34_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_34_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_34_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_35 (
    .io_push_valid      (fifoGroup_35_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_35_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_35_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_35_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_35_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_35_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_35_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_35_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_36 (
    .io_push_valid      (fifoGroup_36_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_36_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_36_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_36_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_36_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_36_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_36_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_36_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_37 (
    .io_push_valid      (fifoGroup_37_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_37_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_37_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_37_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_37_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_37_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_37_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_37_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_38 (
    .io_push_valid      (fifoGroup_38_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_38_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_38_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_38_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_38_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_38_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_38_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_38_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_39 (
    .io_push_valid      (fifoGroup_39_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_39_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_39_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_39_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_39_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_39_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_39_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_39_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_40 (
    .io_push_valid      (fifoGroup_40_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_40_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_40_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_40_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_40_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_40_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_40_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_40_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_41 (
    .io_push_valid      (fifoGroup_41_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_41_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_41_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_41_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_41_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_41_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_41_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_41_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_42 (
    .io_push_valid      (fifoGroup_42_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_42_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_42_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_42_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_42_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_42_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_42_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_42_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_43 (
    .io_push_valid      (fifoGroup_43_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_43_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_43_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_43_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_43_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_43_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_43_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_43_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_44 (
    .io_push_valid      (fifoGroup_44_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_44_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_44_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_44_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_44_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_44_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_44_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_44_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_45 (
    .io_push_valid      (fifoGroup_45_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_45_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_45_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_45_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_45_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_45_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_45_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_45_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_46 (
    .io_push_valid      (fifoGroup_46_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_46_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_46_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_46_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_46_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_46_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_46_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_46_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_47 (
    .io_push_valid      (fifoGroup_47_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_47_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_47_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_47_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_47_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_47_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_47_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_47_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_48 (
    .io_push_valid      (fifoGroup_48_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_48_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_48_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_48_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_48_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_48_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_48_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_48_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_49 (
    .io_push_valid      (fifoGroup_49_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_49_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_49_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_49_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_49_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_49_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_49_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_49_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_50 (
    .io_push_valid      (fifoGroup_50_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_50_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_50_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_50_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_50_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_50_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_50_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_50_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_51 (
    .io_push_valid      (fifoGroup_51_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_51_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_51_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_51_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_51_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_51_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_51_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_51_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_52 (
    .io_push_valid      (fifoGroup_52_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_52_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_52_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_52_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_52_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_52_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_52_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_52_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_53 (
    .io_push_valid      (fifoGroup_53_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_53_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_53_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_53_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_53_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_53_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_53_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_53_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_54 (
    .io_push_valid      (fifoGroup_54_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_54_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_54_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_54_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_54_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_54_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_54_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_54_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_55 (
    .io_push_valid      (fifoGroup_55_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_55_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_55_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_55_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_55_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_55_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_55_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_55_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_56 (
    .io_push_valid      (fifoGroup_56_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_56_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_56_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_56_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_56_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_56_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_56_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_56_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_57 (
    .io_push_valid      (fifoGroup_57_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_57_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_57_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_57_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_57_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_57_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_57_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_57_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_58 (
    .io_push_valid      (fifoGroup_58_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_58_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_58_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_58_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_58_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_58_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_58_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_58_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_59 (
    .io_push_valid      (fifoGroup_59_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_59_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_59_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_59_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_59_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_59_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_59_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_59_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_60 (
    .io_push_valid      (fifoGroup_60_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_60_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_60_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_60_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_60_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_60_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_60_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_60_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_61 (
    .io_push_valid      (fifoGroup_61_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_61_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_61_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_61_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_61_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_61_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_61_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_61_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_62 (
    .io_push_valid      (fifoGroup_62_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_62_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_62_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_62_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_62_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_62_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_62_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_62_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  StreamFifo fifoGroup_63 (
    .io_push_valid      (fifoGroup_63_io_push_valid          ), //i
    .io_push_ready      (fifoGroup_63_io_push_ready          ), //o
    .io_push_payload    (fifoGroup_63_io_push_payload[31:0]  ), //i
    .io_pop_valid       (fifoGroup_63_io_pop_valid           ), //o
    .io_pop_ready       (fifoGroup_63_io_pop_ready           ), //i
    .io_pop_payload     (fifoGroup_63_io_pop_payload[31:0]   ), //o
    .io_flush           (1'b0                                ), //i
    .io_occupancy       (fifoGroup_63_io_occupancy[6:0]      ), //o
    .io_availability    (fifoGroup_63_io_availability[6:0]   ), //o
    .clk                (clk                                 ), //i
    .resetn             (resetn                              )  //i
  );
  always @(*) begin
    case(selectWriteFifo)
      6'b000000 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_0_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_0_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_0_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_0_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_0_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_1_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_1_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_1_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_1_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_1_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_2_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_2_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_2_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_2_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_2_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_3_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_3_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_3_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_3_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_3_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_4_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_4_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_4_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_4_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_4_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_5_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_5_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_5_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_5_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_5_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_6_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_6_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_6_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_6_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_6_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_7_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_7_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_7_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_7_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_7_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_8_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_8_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_8_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_8_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_8_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_9_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_9_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_9_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_9_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_9_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_10_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_10_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_10_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_10_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_10_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_11_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_11_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_11_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_11_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_11_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_12_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_12_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_12_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_12_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_12_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_13_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_13_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_13_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_13_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_13_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_14_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_14_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_14_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_14_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_14_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_15_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_15_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_15_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_15_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_15_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_16_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_16_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_16_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_16_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_16_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_17_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_17_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_17_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_17_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_17_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_18_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_18_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_18_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_18_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_18_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_19_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_19_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_19_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_19_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_19_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_20_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_20_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_20_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_20_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_20_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_21_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_21_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_21_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_21_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_21_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_22_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_22_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_22_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_22_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_22_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_23_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_23_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_23_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_23_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_23_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_24_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_24_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_24_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_24_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_24_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_25_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_25_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_25_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_25_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_25_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_26_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_26_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_26_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_26_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_26_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_27_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_27_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_27_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_27_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_27_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_28_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_28_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_28_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_28_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_28_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_29_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_29_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_29_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_29_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_29_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_30_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_30_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_30_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_30_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_30_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_31_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_31_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_31_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_31_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_31_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_32_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_32_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_32_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_32_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_32_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_33_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_33_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_33_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_33_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_33_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_34_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_34_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_34_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_34_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_34_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_35_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_35_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_35_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_35_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_35_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_36_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_36_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_36_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_36_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_36_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_37_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_37_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_37_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_37_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_37_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_38_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_38_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_38_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_38_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_38_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_39_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_39_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_39_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_39_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_39_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_40_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_40_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_40_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_40_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_40_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_41_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_41_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_41_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_41_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_41_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_42_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_42_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_42_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_42_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_42_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_43_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_43_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_43_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_43_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_43_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_44_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_44_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_44_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_44_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_44_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_45_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_45_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_45_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_45_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_45_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_46_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_46_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_46_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_46_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_46_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_47_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_47_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_47_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_47_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_47_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_48_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_48_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_48_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_48_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_48_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_49_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_49_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_49_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_49_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_49_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_50_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_50_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_50_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_50_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_50_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_51_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_51_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_51_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_51_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_51_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_52_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_52_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_52_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_52_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_52_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_53_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_53_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_53_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_53_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_53_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_54_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_54_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_54_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_54_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_54_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_55_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_55_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_55_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_55_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_55_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_56_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_56_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_56_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_56_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_56_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_57_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_57_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_57_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_57_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_57_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_58_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_58_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_58_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_58_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_58_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_59_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_59_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_59_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_59_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_59_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_60_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_60_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_60_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_60_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_60_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_61_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_61_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_61_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_61_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_61_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l211 = fifoGroup_62_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_62_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_62_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_62_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_62_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l211 = fifoGroup_63_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_63_io_push_ready;
        _zz_when_ArraySlice_l215 = fifoGroup_63_io_occupancy;
        _zz_when_ArraySlice_l334 = fifoGroup_63_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_63_io_push_ready;
        _zz_when_ArraySlice_l338 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l374_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l374 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l374 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_0_valid)
      6'b000000 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_0_valid_2 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_0_payload = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l380_3)
      6'b000000 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l380_2 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l389_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l389 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l389 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l409_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l409 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l409 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l374_1_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l374_1_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_1_valid)
      6'b000000 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_1_valid_2 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_1_payload = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l380_1_4)
      6'b000000 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l380_1_3 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l389_1_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l389_1_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l409_1_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l409_1_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l374_2_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l374_2_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_2_valid)
      6'b000000 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_2_valid_2 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_2_payload = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l380_2_4)
      6'b000000 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l380_2_3 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l389_2_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l389_2_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l409_2_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l409_2_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l374_3_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l374_3_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_3_valid)
      6'b000000 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_3_valid_2 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_3_payload = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l380_3_4)
      6'b000000 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l380_3_3 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l389_3_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l389_3_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l409_3_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l409_3_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l374_4_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l374_4 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_4_valid)
      6'b000000 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_4_valid_2 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_4_payload = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l380_4_4)
      6'b000000 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l380_4_3 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l389_4_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l389_4_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l409_4_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l409_4 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l374_5_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l374_5 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_5_valid)
      6'b000000 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_5_valid_2 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_5_payload = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l380_5_4)
      6'b000000 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l380_5_3 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l389_5_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l389_5_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l409_5_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l409_5 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l374_6_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l374_6 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_6_valid)
      6'b000000 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_6_valid_2 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_6_payload = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l380_6_3)
      6'b000000 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l380_6_2 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l389_6_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l389_6 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l409_6_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l409_6 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l374_7_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l374_7 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_7_valid)
      6'b000000 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_7_valid_2 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_7_payload = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l380_7_3)
      6'b000000 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l380_7_2 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l389_7_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l389_7 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l409_7_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l409_7 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l241_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l241 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l241 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_0_valid_1)
      6'b000000 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_0_valid_3 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_0_payload_1 = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l247_3)
      6'b000000 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l247_2 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l256_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l256 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l256 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l276_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l276 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l276 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l241_1_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l241_1_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_1_valid_1)
      6'b000000 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_1_valid_3 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_1_payload_1 = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l247_1_4)
      6'b000000 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l247_1_3 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l256_1_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l256_1_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l276_1_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l276_1_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l241_2_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l241_2_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_2_valid_1)
      6'b000000 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_2_valid_3 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_2_payload_1 = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l247_2_4)
      6'b000000 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l247_2_3 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l256_2_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l256_2_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l276_2_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l276_2_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l241_3_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l241_3_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_3_valid_1)
      6'b000000 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_3_valid_3 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_3_payload_1 = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l247_3_4)
      6'b000000 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l247_3_3 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l256_3_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l256_3_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l276_3_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l276_3_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l241_4_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l241_4 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_4_valid_1)
      6'b000000 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_4_valid_3 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_4_payload_1 = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l247_4_4)
      6'b000000 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l247_4_3 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l256_4_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l256_4_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l276_4_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l276_4 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l241_5_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l241_5 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_5_valid_1)
      6'b000000 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_5_valid_3 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_5_payload_1 = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l247_5_4)
      6'b000000 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l247_5_3 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l256_5_2)
      6'b000000 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l256_5_1 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l276_5_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l276_5 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l241_6_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l241_6 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_6_valid_1)
      6'b000000 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_6_valid_3 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_6_payload_1 = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l247_6_3)
      6'b000000 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l247_6_2 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l256_6_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l256_6 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l276_6_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l276_6 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l241_7_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l241_7 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_7_valid_1)
      6'b000000 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_0_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_0_io_pop_payload;
      end
      6'b000001 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_1_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_1_io_pop_payload;
      end
      6'b000010 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_2_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_2_io_pop_payload;
      end
      6'b000011 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_3_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_3_io_pop_payload;
      end
      6'b000100 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_4_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_4_io_pop_payload;
      end
      6'b000101 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_5_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_5_io_pop_payload;
      end
      6'b000110 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_6_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_6_io_pop_payload;
      end
      6'b000111 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_7_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_7_io_pop_payload;
      end
      6'b001000 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_8_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_8_io_pop_payload;
      end
      6'b001001 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_9_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_9_io_pop_payload;
      end
      6'b001010 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_10_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_10_io_pop_payload;
      end
      6'b001011 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_11_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_11_io_pop_payload;
      end
      6'b001100 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_12_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_12_io_pop_payload;
      end
      6'b001101 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_13_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_13_io_pop_payload;
      end
      6'b001110 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_14_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_14_io_pop_payload;
      end
      6'b001111 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_15_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_15_io_pop_payload;
      end
      6'b010000 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_16_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_16_io_pop_payload;
      end
      6'b010001 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_17_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_17_io_pop_payload;
      end
      6'b010010 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_18_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_18_io_pop_payload;
      end
      6'b010011 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_19_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_19_io_pop_payload;
      end
      6'b010100 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_20_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_20_io_pop_payload;
      end
      6'b010101 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_21_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_21_io_pop_payload;
      end
      6'b010110 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_22_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_22_io_pop_payload;
      end
      6'b010111 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_23_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_23_io_pop_payload;
      end
      6'b011000 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_24_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_24_io_pop_payload;
      end
      6'b011001 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_25_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_25_io_pop_payload;
      end
      6'b011010 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_26_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_26_io_pop_payload;
      end
      6'b011011 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_27_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_27_io_pop_payload;
      end
      6'b011100 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_28_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_28_io_pop_payload;
      end
      6'b011101 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_29_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_29_io_pop_payload;
      end
      6'b011110 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_30_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_30_io_pop_payload;
      end
      6'b011111 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_31_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_31_io_pop_payload;
      end
      6'b100000 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_32_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_32_io_pop_payload;
      end
      6'b100001 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_33_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_33_io_pop_payload;
      end
      6'b100010 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_34_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_34_io_pop_payload;
      end
      6'b100011 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_35_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_35_io_pop_payload;
      end
      6'b100100 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_36_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_36_io_pop_payload;
      end
      6'b100101 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_37_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_37_io_pop_payload;
      end
      6'b100110 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_38_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_38_io_pop_payload;
      end
      6'b100111 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_39_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_39_io_pop_payload;
      end
      6'b101000 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_40_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_40_io_pop_payload;
      end
      6'b101001 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_41_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_41_io_pop_payload;
      end
      6'b101010 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_42_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_42_io_pop_payload;
      end
      6'b101011 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_43_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_43_io_pop_payload;
      end
      6'b101100 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_44_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_44_io_pop_payload;
      end
      6'b101101 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_45_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_45_io_pop_payload;
      end
      6'b101110 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_46_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_46_io_pop_payload;
      end
      6'b101111 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_47_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_47_io_pop_payload;
      end
      6'b110000 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_48_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_48_io_pop_payload;
      end
      6'b110001 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_49_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_49_io_pop_payload;
      end
      6'b110010 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_50_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_50_io_pop_payload;
      end
      6'b110011 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_51_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_51_io_pop_payload;
      end
      6'b110100 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_52_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_52_io_pop_payload;
      end
      6'b110101 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_53_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_53_io_pop_payload;
      end
      6'b110110 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_54_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_54_io_pop_payload;
      end
      6'b110111 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_55_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_55_io_pop_payload;
      end
      6'b111000 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_56_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_56_io_pop_payload;
      end
      6'b111001 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_57_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_57_io_pop_payload;
      end
      6'b111010 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_58_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_58_io_pop_payload;
      end
      6'b111011 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_59_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_59_io_pop_payload;
      end
      6'b111100 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_60_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_60_io_pop_payload;
      end
      6'b111101 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_61_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_61_io_pop_payload;
      end
      6'b111110 : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_62_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_62_io_pop_payload;
      end
      default : begin
        _zz_outputStreamArrayData_7_valid_3 = fifoGroup_63_io_pop_valid;
        _zz_outputStreamArrayData_7_payload_1 = fifoGroup_63_io_pop_payload;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l247_7_3)
      6'b000000 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l247_7_2 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l256_7_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l256_7 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l276_7_1)
      6'b000000 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_0_io_occupancy;
      end
      6'b000001 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_1_io_occupancy;
      end
      6'b000010 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_2_io_occupancy;
      end
      6'b000011 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_3_io_occupancy;
      end
      6'b000100 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_4_io_occupancy;
      end
      6'b000101 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_5_io_occupancy;
      end
      6'b000110 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_6_io_occupancy;
      end
      6'b000111 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_7_io_occupancy;
      end
      6'b001000 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_8_io_occupancy;
      end
      6'b001001 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_9_io_occupancy;
      end
      6'b001010 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_10_io_occupancy;
      end
      6'b001011 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_11_io_occupancy;
      end
      6'b001100 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_12_io_occupancy;
      end
      6'b001101 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_13_io_occupancy;
      end
      6'b001110 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_14_io_occupancy;
      end
      6'b001111 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_15_io_occupancy;
      end
      6'b010000 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_16_io_occupancy;
      end
      6'b010001 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_17_io_occupancy;
      end
      6'b010010 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_18_io_occupancy;
      end
      6'b010011 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_19_io_occupancy;
      end
      6'b010100 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_20_io_occupancy;
      end
      6'b010101 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_21_io_occupancy;
      end
      6'b010110 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_22_io_occupancy;
      end
      6'b010111 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_23_io_occupancy;
      end
      6'b011000 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_24_io_occupancy;
      end
      6'b011001 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_25_io_occupancy;
      end
      6'b011010 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_26_io_occupancy;
      end
      6'b011011 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_27_io_occupancy;
      end
      6'b011100 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_28_io_occupancy;
      end
      6'b011101 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_29_io_occupancy;
      end
      6'b011110 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_30_io_occupancy;
      end
      6'b011111 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_31_io_occupancy;
      end
      6'b100000 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_32_io_occupancy;
      end
      6'b100001 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_33_io_occupancy;
      end
      6'b100010 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_34_io_occupancy;
      end
      6'b100011 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_35_io_occupancy;
      end
      6'b100100 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_36_io_occupancy;
      end
      6'b100101 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_37_io_occupancy;
      end
      6'b100110 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_38_io_occupancy;
      end
      6'b100111 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_39_io_occupancy;
      end
      6'b101000 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_40_io_occupancy;
      end
      6'b101001 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_41_io_occupancy;
      end
      6'b101010 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_42_io_occupancy;
      end
      6'b101011 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_43_io_occupancy;
      end
      6'b101100 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_44_io_occupancy;
      end
      6'b101101 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_45_io_occupancy;
      end
      6'b101110 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_46_io_occupancy;
      end
      6'b101111 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_47_io_occupancy;
      end
      6'b110000 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_48_io_occupancy;
      end
      6'b110001 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_49_io_occupancy;
      end
      6'b110010 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_50_io_occupancy;
      end
      6'b110011 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_51_io_occupancy;
      end
      6'b110100 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_52_io_occupancy;
      end
      6'b110101 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_53_io_occupancy;
      end
      6'b110110 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_54_io_occupancy;
      end
      6'b110111 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_55_io_occupancy;
      end
      6'b111000 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_56_io_occupancy;
      end
      6'b111001 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_57_io_occupancy;
      end
      6'b111010 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_58_io_occupancy;
      end
      6'b111011 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_59_io_occupancy;
      end
      6'b111100 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_60_io_occupancy;
      end
      6'b111101 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_61_io_occupancy;
      end
      6'b111110 : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_62_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l276_7 = fifoGroup_63_io_occupancy;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_BOOT : arraySliceStateMachine_stateReg_string = "BOOT         ";
      arraySliceStateMachine_enumDef_writeDataOnly : arraySliceStateMachine_stateReg_string = "writeDataOnly";
      arraySliceStateMachine_enumDef_readDataOnly : arraySliceStateMachine_stateReg_string = "readDataOnly ";
      arraySliceStateMachine_enumDef_readWriteData : arraySliceStateMachine_stateReg_string = "readWriteData";
      default : arraySliceStateMachine_stateReg_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(arraySliceStateMachine_stateNext)
      arraySliceStateMachine_enumDef_BOOT : arraySliceStateMachine_stateNext_string = "BOOT         ";
      arraySliceStateMachine_enumDef_writeDataOnly : arraySliceStateMachine_stateNext_string = "writeDataOnly";
      arraySliceStateMachine_enumDef_readDataOnly : arraySliceStateMachine_stateNext_string = "readDataOnly ";
      arraySliceStateMachine_enumDef_readWriteData : arraySliceStateMachine_stateNext_string = "readWriteData";
      default : arraySliceStateMachine_stateNext_string = "?????????????";
    endcase
  end
  `endif

  always @(*) begin
    handshakeTimes_0_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_0_fire_6) begin
          if(!when_ArraySlice_l455) begin
            handshakeTimes_0_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_0_fire_13) begin
          if(!when_ArraySlice_l322) begin
            handshakeTimes_0_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_0_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_0_fire_6) begin
          if(when_ArraySlice_l455) begin
            handshakeTimes_0_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_0_fire_13) begin
          if(when_ArraySlice_l322) begin
            handshakeTimes_0_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_0_willOverflowIfInc = (handshakeTimes_0_value == 13'h1000);
  assign handshakeTimes_0_willOverflow = (handshakeTimes_0_willOverflowIfInc && handshakeTimes_0_willIncrement);
  always @(*) begin
    if(handshakeTimes_0_willOverflow) begin
      handshakeTimes_0_valueNext = 13'h0;
    end else begin
      handshakeTimes_0_valueNext = (handshakeTimes_0_value + _zz_handshakeTimes_0_valueNext);
    end
    if(handshakeTimes_0_willClear) begin
      handshakeTimes_0_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_1_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_1_fire_6) begin
          if(!when_ArraySlice_l455_1) begin
            handshakeTimes_1_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_1_fire_13) begin
          if(!when_ArraySlice_l322_1) begin
            handshakeTimes_1_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_1_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_1_fire_6) begin
          if(when_ArraySlice_l455_1) begin
            handshakeTimes_1_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_1_fire_13) begin
          if(when_ArraySlice_l322_1) begin
            handshakeTimes_1_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_1_willOverflowIfInc = (handshakeTimes_1_value == 13'h1000);
  assign handshakeTimes_1_willOverflow = (handshakeTimes_1_willOverflowIfInc && handshakeTimes_1_willIncrement);
  always @(*) begin
    if(handshakeTimes_1_willOverflow) begin
      handshakeTimes_1_valueNext = 13'h0;
    end else begin
      handshakeTimes_1_valueNext = (handshakeTimes_1_value + _zz_handshakeTimes_1_valueNext);
    end
    if(handshakeTimes_1_willClear) begin
      handshakeTimes_1_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_2_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_2_fire_6) begin
          if(!when_ArraySlice_l455_2) begin
            handshakeTimes_2_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_2_fire_13) begin
          if(!when_ArraySlice_l322_2) begin
            handshakeTimes_2_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_2_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_2_fire_6) begin
          if(when_ArraySlice_l455_2) begin
            handshakeTimes_2_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_2_fire_13) begin
          if(when_ArraySlice_l322_2) begin
            handshakeTimes_2_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_2_willOverflowIfInc = (handshakeTimes_2_value == 13'h1000);
  assign handshakeTimes_2_willOverflow = (handshakeTimes_2_willOverflowIfInc && handshakeTimes_2_willIncrement);
  always @(*) begin
    if(handshakeTimes_2_willOverflow) begin
      handshakeTimes_2_valueNext = 13'h0;
    end else begin
      handshakeTimes_2_valueNext = (handshakeTimes_2_value + _zz_handshakeTimes_2_valueNext);
    end
    if(handshakeTimes_2_willClear) begin
      handshakeTimes_2_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_3_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_3_fire_6) begin
          if(!when_ArraySlice_l455_3) begin
            handshakeTimes_3_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_3_fire_13) begin
          if(!when_ArraySlice_l322_3) begin
            handshakeTimes_3_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_3_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_3_fire_6) begin
          if(when_ArraySlice_l455_3) begin
            handshakeTimes_3_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_3_fire_13) begin
          if(when_ArraySlice_l322_3) begin
            handshakeTimes_3_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_3_willOverflowIfInc = (handshakeTimes_3_value == 13'h1000);
  assign handshakeTimes_3_willOverflow = (handshakeTimes_3_willOverflowIfInc && handshakeTimes_3_willIncrement);
  always @(*) begin
    if(handshakeTimes_3_willOverflow) begin
      handshakeTimes_3_valueNext = 13'h0;
    end else begin
      handshakeTimes_3_valueNext = (handshakeTimes_3_value + _zz_handshakeTimes_3_valueNext);
    end
    if(handshakeTimes_3_willClear) begin
      handshakeTimes_3_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_4_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_4_fire_6) begin
          if(!when_ArraySlice_l455_4) begin
            handshakeTimes_4_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_4_fire_13) begin
          if(!when_ArraySlice_l322_4) begin
            handshakeTimes_4_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_4_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_4_fire_6) begin
          if(when_ArraySlice_l455_4) begin
            handshakeTimes_4_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_4_fire_13) begin
          if(when_ArraySlice_l322_4) begin
            handshakeTimes_4_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_4_willOverflowIfInc = (handshakeTimes_4_value == 13'h1000);
  assign handshakeTimes_4_willOverflow = (handshakeTimes_4_willOverflowIfInc && handshakeTimes_4_willIncrement);
  always @(*) begin
    if(handshakeTimes_4_willOverflow) begin
      handshakeTimes_4_valueNext = 13'h0;
    end else begin
      handshakeTimes_4_valueNext = (handshakeTimes_4_value + _zz_handshakeTimes_4_valueNext);
    end
    if(handshakeTimes_4_willClear) begin
      handshakeTimes_4_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_5_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_5_fire_6) begin
          if(!when_ArraySlice_l455_5) begin
            handshakeTimes_5_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_5_fire_13) begin
          if(!when_ArraySlice_l322_5) begin
            handshakeTimes_5_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_5_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_5_fire_6) begin
          if(when_ArraySlice_l455_5) begin
            handshakeTimes_5_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_5_fire_13) begin
          if(when_ArraySlice_l322_5) begin
            handshakeTimes_5_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_5_willOverflowIfInc = (handshakeTimes_5_value == 13'h1000);
  assign handshakeTimes_5_willOverflow = (handshakeTimes_5_willOverflowIfInc && handshakeTimes_5_willIncrement);
  always @(*) begin
    if(handshakeTimes_5_willOverflow) begin
      handshakeTimes_5_valueNext = 13'h0;
    end else begin
      handshakeTimes_5_valueNext = (handshakeTimes_5_value + _zz_handshakeTimes_5_valueNext);
    end
    if(handshakeTimes_5_willClear) begin
      handshakeTimes_5_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_6_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_6_fire_6) begin
          if(!when_ArraySlice_l455_6) begin
            handshakeTimes_6_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_6_fire_13) begin
          if(!when_ArraySlice_l322_6) begin
            handshakeTimes_6_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_6_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_6_fire_6) begin
          if(when_ArraySlice_l455_6) begin
            handshakeTimes_6_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_6_fire_13) begin
          if(when_ArraySlice_l322_6) begin
            handshakeTimes_6_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_6_willOverflowIfInc = (handshakeTimes_6_value == 13'h1000);
  assign handshakeTimes_6_willOverflow = (handshakeTimes_6_willOverflowIfInc && handshakeTimes_6_willIncrement);
  always @(*) begin
    if(handshakeTimes_6_willOverflow) begin
      handshakeTimes_6_valueNext = 13'h0;
    end else begin
      handshakeTimes_6_valueNext = (handshakeTimes_6_value + _zz_handshakeTimes_6_valueNext);
    end
    if(handshakeTimes_6_willClear) begin
      handshakeTimes_6_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_7_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_7_fire_6) begin
          if(!when_ArraySlice_l455_7) begin
            handshakeTimes_7_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_7_fire_13) begin
          if(!when_ArraySlice_l322_7) begin
            handshakeTimes_7_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_7_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_7_fire_6) begin
          if(when_ArraySlice_l455_7) begin
            handshakeTimes_7_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_7_fire_13) begin
          if(when_ArraySlice_l322_7) begin
            handshakeTimes_7_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_7_willOverflowIfInc = (handshakeTimes_7_value == 13'h1000);
  assign handshakeTimes_7_willOverflow = (handshakeTimes_7_willOverflowIfInc && handshakeTimes_7_willIncrement);
  always @(*) begin
    if(handshakeTimes_7_willOverflow) begin
      handshakeTimes_7_valueNext = 13'h0;
    end else begin
      handshakeTimes_7_valueNext = (handshakeTimes_7_value + _zz_handshakeTimes_7_valueNext);
    end
    if(handshakeTimes_7_willClear) begin
      handshakeTimes_7_valueNext = 13'h0;
    end
  end

  always @(*) begin
    outSliceNumb_0_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l379) begin
            if(when_ArraySlice_l380) begin
              if(when_ArraySlice_l381) begin
                outSliceNumb_0_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l389) begin
              if(when_ArraySlice_l390) begin
                if(when_ArraySlice_l392) begin
                  outSliceNumb_0_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409) begin
              if(when_ArraySlice_l410) begin
                if(when_ArraySlice_l412) begin
                  outSliceNumb_0_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434) begin
            if(when_ArraySlice_l436) begin
              if(when_ArraySlice_l437) begin
                outSliceNumb_0_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l246) begin
            if(when_ArraySlice_l247) begin
              if(when_ArraySlice_l248) begin
                outSliceNumb_0_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l256) begin
              if(when_ArraySlice_l257) begin
                if(when_ArraySlice_l259) begin
                  outSliceNumb_0_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276) begin
              if(when_ArraySlice_l277) begin
                if(when_ArraySlice_l279) begin
                  outSliceNumb_0_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301) begin
            if(when_ArraySlice_l303) begin
              if(when_ArraySlice_l304) begin
                outSliceNumb_0_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_0_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l379) begin
            if(when_ArraySlice_l389) begin
              if(when_ArraySlice_l390) begin
                if(!when_ArraySlice_l392) begin
                  outSliceNumb_0_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409) begin
              if(when_ArraySlice_l410) begin
                if(!when_ArraySlice_l412) begin
                  outSliceNumb_0_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434) begin
            if(when_ArraySlice_l436) begin
              if(!when_ArraySlice_l437) begin
                outSliceNumb_0_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l246) begin
            if(when_ArraySlice_l256) begin
              if(when_ArraySlice_l257) begin
                if(!when_ArraySlice_l259) begin
                  outSliceNumb_0_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276) begin
              if(when_ArraySlice_l277) begin
                if(!when_ArraySlice_l279) begin
                  outSliceNumb_0_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301) begin
            if(when_ArraySlice_l303) begin
              if(!when_ArraySlice_l304) begin
                outSliceNumb_0_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_0_willOverflowIfInc = (outSliceNumb_0_value == 7'h40);
  assign outSliceNumb_0_willOverflow = (outSliceNumb_0_willOverflowIfInc && outSliceNumb_0_willIncrement);
  always @(*) begin
    if(outSliceNumb_0_willOverflow) begin
      outSliceNumb_0_valueNext = 7'h0;
    end else begin
      outSliceNumb_0_valueNext = (outSliceNumb_0_value + _zz_outSliceNumb_0_valueNext);
    end
    if(outSliceNumb_0_willClear) begin
      outSliceNumb_0_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_1_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l379_1) begin
            if(when_ArraySlice_l380_1) begin
              if(when_ArraySlice_l381_1) begin
                outSliceNumb_1_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l389_1) begin
              if(when_ArraySlice_l390_1) begin
                if(when_ArraySlice_l392_1) begin
                  outSliceNumb_1_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_1) begin
              if(when_ArraySlice_l410_1) begin
                if(when_ArraySlice_l412_1) begin
                  outSliceNumb_1_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_1) begin
            if(when_ArraySlice_l436_1) begin
              if(when_ArraySlice_l437_1) begin
                outSliceNumb_1_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l246_1) begin
            if(when_ArraySlice_l247_1) begin
              if(when_ArraySlice_l248_1) begin
                outSliceNumb_1_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l256_1) begin
              if(when_ArraySlice_l257_1) begin
                if(when_ArraySlice_l259_1) begin
                  outSliceNumb_1_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_1) begin
              if(when_ArraySlice_l277_1) begin
                if(when_ArraySlice_l279_1) begin
                  outSliceNumb_1_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_1) begin
            if(when_ArraySlice_l303_1) begin
              if(when_ArraySlice_l304_1) begin
                outSliceNumb_1_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_1_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l379_1) begin
            if(when_ArraySlice_l389_1) begin
              if(when_ArraySlice_l390_1) begin
                if(!when_ArraySlice_l392_1) begin
                  outSliceNumb_1_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_1) begin
              if(when_ArraySlice_l410_1) begin
                if(!when_ArraySlice_l412_1) begin
                  outSliceNumb_1_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_1) begin
            if(when_ArraySlice_l436_1) begin
              if(!when_ArraySlice_l437_1) begin
                outSliceNumb_1_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l246_1) begin
            if(when_ArraySlice_l256_1) begin
              if(when_ArraySlice_l257_1) begin
                if(!when_ArraySlice_l259_1) begin
                  outSliceNumb_1_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_1) begin
              if(when_ArraySlice_l277_1) begin
                if(!when_ArraySlice_l279_1) begin
                  outSliceNumb_1_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_1) begin
            if(when_ArraySlice_l303_1) begin
              if(!when_ArraySlice_l304_1) begin
                outSliceNumb_1_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_1_willOverflowIfInc = (outSliceNumb_1_value == 7'h40);
  assign outSliceNumb_1_willOverflow = (outSliceNumb_1_willOverflowIfInc && outSliceNumb_1_willIncrement);
  always @(*) begin
    if(outSliceNumb_1_willOverflow) begin
      outSliceNumb_1_valueNext = 7'h0;
    end else begin
      outSliceNumb_1_valueNext = (outSliceNumb_1_value + _zz_outSliceNumb_1_valueNext);
    end
    if(outSliceNumb_1_willClear) begin
      outSliceNumb_1_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_2_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l379_2) begin
            if(when_ArraySlice_l380_2) begin
              if(when_ArraySlice_l381_2) begin
                outSliceNumb_2_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l389_2) begin
              if(when_ArraySlice_l390_2) begin
                if(when_ArraySlice_l392_2) begin
                  outSliceNumb_2_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_2) begin
              if(when_ArraySlice_l410_2) begin
                if(when_ArraySlice_l412_2) begin
                  outSliceNumb_2_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_2) begin
            if(when_ArraySlice_l436_2) begin
              if(when_ArraySlice_l437_2) begin
                outSliceNumb_2_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l246_2) begin
            if(when_ArraySlice_l247_2) begin
              if(when_ArraySlice_l248_2) begin
                outSliceNumb_2_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l256_2) begin
              if(when_ArraySlice_l257_2) begin
                if(when_ArraySlice_l259_2) begin
                  outSliceNumb_2_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_2) begin
              if(when_ArraySlice_l277_2) begin
                if(when_ArraySlice_l279_2) begin
                  outSliceNumb_2_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_2) begin
            if(when_ArraySlice_l303_2) begin
              if(when_ArraySlice_l304_2) begin
                outSliceNumb_2_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_2_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l379_2) begin
            if(when_ArraySlice_l389_2) begin
              if(when_ArraySlice_l390_2) begin
                if(!when_ArraySlice_l392_2) begin
                  outSliceNumb_2_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_2) begin
              if(when_ArraySlice_l410_2) begin
                if(!when_ArraySlice_l412_2) begin
                  outSliceNumb_2_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_2) begin
            if(when_ArraySlice_l436_2) begin
              if(!when_ArraySlice_l437_2) begin
                outSliceNumb_2_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l246_2) begin
            if(when_ArraySlice_l256_2) begin
              if(when_ArraySlice_l257_2) begin
                if(!when_ArraySlice_l259_2) begin
                  outSliceNumb_2_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_2) begin
              if(when_ArraySlice_l277_2) begin
                if(!when_ArraySlice_l279_2) begin
                  outSliceNumb_2_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_2) begin
            if(when_ArraySlice_l303_2) begin
              if(!when_ArraySlice_l304_2) begin
                outSliceNumb_2_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_2_willOverflowIfInc = (outSliceNumb_2_value == 7'h40);
  assign outSliceNumb_2_willOverflow = (outSliceNumb_2_willOverflowIfInc && outSliceNumb_2_willIncrement);
  always @(*) begin
    if(outSliceNumb_2_willOverflow) begin
      outSliceNumb_2_valueNext = 7'h0;
    end else begin
      outSliceNumb_2_valueNext = (outSliceNumb_2_value + _zz_outSliceNumb_2_valueNext);
    end
    if(outSliceNumb_2_willClear) begin
      outSliceNumb_2_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_3_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l379_3) begin
            if(when_ArraySlice_l380_3) begin
              if(when_ArraySlice_l381_3) begin
                outSliceNumb_3_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l389_3) begin
              if(when_ArraySlice_l390_3) begin
                if(when_ArraySlice_l392_3) begin
                  outSliceNumb_3_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_3) begin
              if(when_ArraySlice_l410_3) begin
                if(when_ArraySlice_l412_3) begin
                  outSliceNumb_3_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_3) begin
            if(when_ArraySlice_l436_3) begin
              if(when_ArraySlice_l437_3) begin
                outSliceNumb_3_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l246_3) begin
            if(when_ArraySlice_l247_3) begin
              if(when_ArraySlice_l248_3) begin
                outSliceNumb_3_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l256_3) begin
              if(when_ArraySlice_l257_3) begin
                if(when_ArraySlice_l259_3) begin
                  outSliceNumb_3_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_3) begin
              if(when_ArraySlice_l277_3) begin
                if(when_ArraySlice_l279_3) begin
                  outSliceNumb_3_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_3) begin
            if(when_ArraySlice_l303_3) begin
              if(when_ArraySlice_l304_3) begin
                outSliceNumb_3_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_3_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l379_3) begin
            if(when_ArraySlice_l389_3) begin
              if(when_ArraySlice_l390_3) begin
                if(!when_ArraySlice_l392_3) begin
                  outSliceNumb_3_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_3) begin
              if(when_ArraySlice_l410_3) begin
                if(!when_ArraySlice_l412_3) begin
                  outSliceNumb_3_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_3) begin
            if(when_ArraySlice_l436_3) begin
              if(!when_ArraySlice_l437_3) begin
                outSliceNumb_3_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l246_3) begin
            if(when_ArraySlice_l256_3) begin
              if(when_ArraySlice_l257_3) begin
                if(!when_ArraySlice_l259_3) begin
                  outSliceNumb_3_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_3) begin
              if(when_ArraySlice_l277_3) begin
                if(!when_ArraySlice_l279_3) begin
                  outSliceNumb_3_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_3) begin
            if(when_ArraySlice_l303_3) begin
              if(!when_ArraySlice_l304_3) begin
                outSliceNumb_3_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_3_willOverflowIfInc = (outSliceNumb_3_value == 7'h40);
  assign outSliceNumb_3_willOverflow = (outSliceNumb_3_willOverflowIfInc && outSliceNumb_3_willIncrement);
  always @(*) begin
    if(outSliceNumb_3_willOverflow) begin
      outSliceNumb_3_valueNext = 7'h0;
    end else begin
      outSliceNumb_3_valueNext = (outSliceNumb_3_value + _zz_outSliceNumb_3_valueNext);
    end
    if(outSliceNumb_3_willClear) begin
      outSliceNumb_3_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_4_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l379_4) begin
            if(when_ArraySlice_l380_4) begin
              if(when_ArraySlice_l381_4) begin
                outSliceNumb_4_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l389_4) begin
              if(when_ArraySlice_l390_4) begin
                if(when_ArraySlice_l392_4) begin
                  outSliceNumb_4_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_4) begin
              if(when_ArraySlice_l410_4) begin
                if(when_ArraySlice_l412_4) begin
                  outSliceNumb_4_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_4) begin
            if(when_ArraySlice_l436_4) begin
              if(when_ArraySlice_l437_4) begin
                outSliceNumb_4_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l246_4) begin
            if(when_ArraySlice_l247_4) begin
              if(when_ArraySlice_l248_4) begin
                outSliceNumb_4_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l256_4) begin
              if(when_ArraySlice_l257_4) begin
                if(when_ArraySlice_l259_4) begin
                  outSliceNumb_4_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_4) begin
              if(when_ArraySlice_l277_4) begin
                if(when_ArraySlice_l279_4) begin
                  outSliceNumb_4_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_4) begin
            if(when_ArraySlice_l303_4) begin
              if(when_ArraySlice_l304_4) begin
                outSliceNumb_4_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_4_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l379_4) begin
            if(when_ArraySlice_l389_4) begin
              if(when_ArraySlice_l390_4) begin
                if(!when_ArraySlice_l392_4) begin
                  outSliceNumb_4_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_4) begin
              if(when_ArraySlice_l410_4) begin
                if(!when_ArraySlice_l412_4) begin
                  outSliceNumb_4_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_4) begin
            if(when_ArraySlice_l436_4) begin
              if(!when_ArraySlice_l437_4) begin
                outSliceNumb_4_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l246_4) begin
            if(when_ArraySlice_l256_4) begin
              if(when_ArraySlice_l257_4) begin
                if(!when_ArraySlice_l259_4) begin
                  outSliceNumb_4_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_4) begin
              if(when_ArraySlice_l277_4) begin
                if(!when_ArraySlice_l279_4) begin
                  outSliceNumb_4_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_4) begin
            if(when_ArraySlice_l303_4) begin
              if(!when_ArraySlice_l304_4) begin
                outSliceNumb_4_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_4_willOverflowIfInc = (outSliceNumb_4_value == 7'h40);
  assign outSliceNumb_4_willOverflow = (outSliceNumb_4_willOverflowIfInc && outSliceNumb_4_willIncrement);
  always @(*) begin
    if(outSliceNumb_4_willOverflow) begin
      outSliceNumb_4_valueNext = 7'h0;
    end else begin
      outSliceNumb_4_valueNext = (outSliceNumb_4_value + _zz_outSliceNumb_4_valueNext);
    end
    if(outSliceNumb_4_willClear) begin
      outSliceNumb_4_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_5_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l379_5) begin
            if(when_ArraySlice_l380_5) begin
              if(when_ArraySlice_l381_5) begin
                outSliceNumb_5_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l389_5) begin
              if(when_ArraySlice_l390_5) begin
                if(when_ArraySlice_l392_5) begin
                  outSliceNumb_5_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_5) begin
              if(when_ArraySlice_l410_5) begin
                if(when_ArraySlice_l412_5) begin
                  outSliceNumb_5_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_5) begin
            if(when_ArraySlice_l436_5) begin
              if(when_ArraySlice_l437_5) begin
                outSliceNumb_5_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l246_5) begin
            if(when_ArraySlice_l247_5) begin
              if(when_ArraySlice_l248_5) begin
                outSliceNumb_5_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l256_5) begin
              if(when_ArraySlice_l257_5) begin
                if(when_ArraySlice_l259_5) begin
                  outSliceNumb_5_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_5) begin
              if(when_ArraySlice_l277_5) begin
                if(when_ArraySlice_l279_5) begin
                  outSliceNumb_5_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_5) begin
            if(when_ArraySlice_l303_5) begin
              if(when_ArraySlice_l304_5) begin
                outSliceNumb_5_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_5_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l379_5) begin
            if(when_ArraySlice_l389_5) begin
              if(when_ArraySlice_l390_5) begin
                if(!when_ArraySlice_l392_5) begin
                  outSliceNumb_5_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_5) begin
              if(when_ArraySlice_l410_5) begin
                if(!when_ArraySlice_l412_5) begin
                  outSliceNumb_5_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_5) begin
            if(when_ArraySlice_l436_5) begin
              if(!when_ArraySlice_l437_5) begin
                outSliceNumb_5_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l246_5) begin
            if(when_ArraySlice_l256_5) begin
              if(when_ArraySlice_l257_5) begin
                if(!when_ArraySlice_l259_5) begin
                  outSliceNumb_5_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_5) begin
              if(when_ArraySlice_l277_5) begin
                if(!when_ArraySlice_l279_5) begin
                  outSliceNumb_5_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_5) begin
            if(when_ArraySlice_l303_5) begin
              if(!when_ArraySlice_l304_5) begin
                outSliceNumb_5_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_5_willOverflowIfInc = (outSliceNumb_5_value == 7'h40);
  assign outSliceNumb_5_willOverflow = (outSliceNumb_5_willOverflowIfInc && outSliceNumb_5_willIncrement);
  always @(*) begin
    if(outSliceNumb_5_willOverflow) begin
      outSliceNumb_5_valueNext = 7'h0;
    end else begin
      outSliceNumb_5_valueNext = (outSliceNumb_5_value + _zz_outSliceNumb_5_valueNext);
    end
    if(outSliceNumb_5_willClear) begin
      outSliceNumb_5_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_6_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l379_6) begin
            if(when_ArraySlice_l380_6) begin
              if(when_ArraySlice_l381_6) begin
                outSliceNumb_6_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l389_6) begin
              if(when_ArraySlice_l390_6) begin
                if(when_ArraySlice_l392_6) begin
                  outSliceNumb_6_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_6) begin
              if(when_ArraySlice_l410_6) begin
                if(when_ArraySlice_l412_6) begin
                  outSliceNumb_6_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_6) begin
            if(when_ArraySlice_l436_6) begin
              if(when_ArraySlice_l437_6) begin
                outSliceNumb_6_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l246_6) begin
            if(when_ArraySlice_l247_6) begin
              if(when_ArraySlice_l248_6) begin
                outSliceNumb_6_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l256_6) begin
              if(when_ArraySlice_l257_6) begin
                if(when_ArraySlice_l259_6) begin
                  outSliceNumb_6_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_6) begin
              if(when_ArraySlice_l277_6) begin
                if(when_ArraySlice_l279_6) begin
                  outSliceNumb_6_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_6) begin
            if(when_ArraySlice_l303_6) begin
              if(when_ArraySlice_l304_6) begin
                outSliceNumb_6_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_6_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l379_6) begin
            if(when_ArraySlice_l389_6) begin
              if(when_ArraySlice_l390_6) begin
                if(!when_ArraySlice_l392_6) begin
                  outSliceNumb_6_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_6) begin
              if(when_ArraySlice_l410_6) begin
                if(!when_ArraySlice_l412_6) begin
                  outSliceNumb_6_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_6) begin
            if(when_ArraySlice_l436_6) begin
              if(!when_ArraySlice_l437_6) begin
                outSliceNumb_6_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l246_6) begin
            if(when_ArraySlice_l256_6) begin
              if(when_ArraySlice_l257_6) begin
                if(!when_ArraySlice_l259_6) begin
                  outSliceNumb_6_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_6) begin
              if(when_ArraySlice_l277_6) begin
                if(!when_ArraySlice_l279_6) begin
                  outSliceNumb_6_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_6) begin
            if(when_ArraySlice_l303_6) begin
              if(!when_ArraySlice_l304_6) begin
                outSliceNumb_6_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_6_willOverflowIfInc = (outSliceNumb_6_value == 7'h40);
  assign outSliceNumb_6_willOverflow = (outSliceNumb_6_willOverflowIfInc && outSliceNumb_6_willIncrement);
  always @(*) begin
    if(outSliceNumb_6_willOverflow) begin
      outSliceNumb_6_valueNext = 7'h0;
    end else begin
      outSliceNumb_6_valueNext = (outSliceNumb_6_value + _zz_outSliceNumb_6_valueNext);
    end
    if(outSliceNumb_6_willClear) begin
      outSliceNumb_6_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_7_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l379_7) begin
            if(when_ArraySlice_l380_7) begin
              if(when_ArraySlice_l381_7) begin
                outSliceNumb_7_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l389_7) begin
              if(when_ArraySlice_l390_7) begin
                if(when_ArraySlice_l392_7) begin
                  outSliceNumb_7_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_7) begin
              if(when_ArraySlice_l410_7) begin
                if(when_ArraySlice_l412_7) begin
                  outSliceNumb_7_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_7) begin
            if(when_ArraySlice_l436_7) begin
              if(when_ArraySlice_l437_7) begin
                outSliceNumb_7_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l246_7) begin
            if(when_ArraySlice_l247_7) begin
              if(when_ArraySlice_l248_7) begin
                outSliceNumb_7_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l256_7) begin
              if(when_ArraySlice_l257_7) begin
                if(when_ArraySlice_l259_7) begin
                  outSliceNumb_7_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_7) begin
              if(when_ArraySlice_l277_7) begin
                if(when_ArraySlice_l279_7) begin
                  outSliceNumb_7_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_7) begin
            if(when_ArraySlice_l303_7) begin
              if(when_ArraySlice_l304_7) begin
                outSliceNumb_7_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_7_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l379_7) begin
            if(when_ArraySlice_l389_7) begin
              if(when_ArraySlice_l390_7) begin
                if(!when_ArraySlice_l392_7) begin
                  outSliceNumb_7_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l409_7) begin
              if(when_ArraySlice_l410_7) begin
                if(!when_ArraySlice_l412_7) begin
                  outSliceNumb_7_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l434_7) begin
            if(when_ArraySlice_l436_7) begin
              if(!when_ArraySlice_l437_7) begin
                outSliceNumb_7_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l246_7) begin
            if(when_ArraySlice_l256_7) begin
              if(when_ArraySlice_l257_7) begin
                if(!when_ArraySlice_l259_7) begin
                  outSliceNumb_7_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l276_7) begin
              if(when_ArraySlice_l277_7) begin
                if(!when_ArraySlice_l279_7) begin
                  outSliceNumb_7_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l301_7) begin
            if(when_ArraySlice_l303_7) begin
              if(!when_ArraySlice_l304_7) begin
                outSliceNumb_7_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_7_willOverflowIfInc = (outSliceNumb_7_value == 7'h40);
  assign outSliceNumb_7_willOverflow = (outSliceNumb_7_willOverflowIfInc && outSliceNumb_7_willIncrement);
  always @(*) begin
    if(outSliceNumb_7_willOverflow) begin
      outSliceNumb_7_valueNext = 7'h0;
    end else begin
      outSliceNumb_7_valueNext = (outSliceNumb_7_value + _zz_outSliceNumb_7_valueNext);
    end
    if(outSliceNumb_7_willClear) begin
      outSliceNumb_7_valueNext = 7'h0;
    end
  end

  always @(*) begin
    inputStreamArrayData_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          inputStreamArrayData_ready = _zz_inputStreamArrayData_ready;
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            inputStreamArrayData_ready = _zz_inputStreamArrayData_ready_1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_0_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            outputStreamArrayData_0_valid = _zz_outputStreamArrayData_0_valid_2;
          end
          if(when_ArraySlice_l379) begin
            if(when_ArraySlice_l409) begin
              outputStreamArrayData_0_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l434) begin
            outputStreamArrayData_0_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            outputStreamArrayData_0_valid = _zz_outputStreamArrayData_0_valid_3;
          end
          if(when_ArraySlice_l246) begin
            if(when_ArraySlice_l276) begin
              outputStreamArrayData_0_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l301) begin
            outputStreamArrayData_0_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_0_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            outputStreamArrayData_0_payload = _zz_outputStreamArrayData_0_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            outputStreamArrayData_0_payload = _zz_outputStreamArrayData_0_payload_1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_1_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            outputStreamArrayData_1_valid = _zz_outputStreamArrayData_1_valid_2;
          end
          if(when_ArraySlice_l379_1) begin
            if(when_ArraySlice_l409_1) begin
              outputStreamArrayData_1_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l434_1) begin
            outputStreamArrayData_1_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            outputStreamArrayData_1_valid = _zz_outputStreamArrayData_1_valid_3;
          end
          if(when_ArraySlice_l246_1) begin
            if(when_ArraySlice_l276_1) begin
              outputStreamArrayData_1_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l301_1) begin
            outputStreamArrayData_1_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_1_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            outputStreamArrayData_1_payload = _zz_outputStreamArrayData_1_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            outputStreamArrayData_1_payload = _zz_outputStreamArrayData_1_payload_1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_2_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            outputStreamArrayData_2_valid = _zz_outputStreamArrayData_2_valid_2;
          end
          if(when_ArraySlice_l379_2) begin
            if(when_ArraySlice_l409_2) begin
              outputStreamArrayData_2_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l434_2) begin
            outputStreamArrayData_2_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            outputStreamArrayData_2_valid = _zz_outputStreamArrayData_2_valid_3;
          end
          if(when_ArraySlice_l246_2) begin
            if(when_ArraySlice_l276_2) begin
              outputStreamArrayData_2_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l301_2) begin
            outputStreamArrayData_2_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_2_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            outputStreamArrayData_2_payload = _zz_outputStreamArrayData_2_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            outputStreamArrayData_2_payload = _zz_outputStreamArrayData_2_payload_1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_3_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            outputStreamArrayData_3_valid = _zz_outputStreamArrayData_3_valid_2;
          end
          if(when_ArraySlice_l379_3) begin
            if(when_ArraySlice_l409_3) begin
              outputStreamArrayData_3_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l434_3) begin
            outputStreamArrayData_3_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            outputStreamArrayData_3_valid = _zz_outputStreamArrayData_3_valid_3;
          end
          if(when_ArraySlice_l246_3) begin
            if(when_ArraySlice_l276_3) begin
              outputStreamArrayData_3_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l301_3) begin
            outputStreamArrayData_3_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_3_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            outputStreamArrayData_3_payload = _zz_outputStreamArrayData_3_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            outputStreamArrayData_3_payload = _zz_outputStreamArrayData_3_payload_1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_4_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            outputStreamArrayData_4_valid = _zz_outputStreamArrayData_4_valid_2;
          end
          if(when_ArraySlice_l379_4) begin
            if(when_ArraySlice_l409_4) begin
              outputStreamArrayData_4_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l434_4) begin
            outputStreamArrayData_4_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            outputStreamArrayData_4_valid = _zz_outputStreamArrayData_4_valid_3;
          end
          if(when_ArraySlice_l246_4) begin
            if(when_ArraySlice_l276_4) begin
              outputStreamArrayData_4_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l301_4) begin
            outputStreamArrayData_4_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_4_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            outputStreamArrayData_4_payload = _zz_outputStreamArrayData_4_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            outputStreamArrayData_4_payload = _zz_outputStreamArrayData_4_payload_1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_5_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            outputStreamArrayData_5_valid = _zz_outputStreamArrayData_5_valid_2;
          end
          if(when_ArraySlice_l379_5) begin
            if(when_ArraySlice_l409_5) begin
              outputStreamArrayData_5_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l434_5) begin
            outputStreamArrayData_5_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            outputStreamArrayData_5_valid = _zz_outputStreamArrayData_5_valid_3;
          end
          if(when_ArraySlice_l246_5) begin
            if(when_ArraySlice_l276_5) begin
              outputStreamArrayData_5_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l301_5) begin
            outputStreamArrayData_5_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_5_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            outputStreamArrayData_5_payload = _zz_outputStreamArrayData_5_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            outputStreamArrayData_5_payload = _zz_outputStreamArrayData_5_payload_1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_6_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            outputStreamArrayData_6_valid = _zz_outputStreamArrayData_6_valid_2;
          end
          if(when_ArraySlice_l379_6) begin
            if(when_ArraySlice_l409_6) begin
              outputStreamArrayData_6_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l434_6) begin
            outputStreamArrayData_6_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            outputStreamArrayData_6_valid = _zz_outputStreamArrayData_6_valid_3;
          end
          if(when_ArraySlice_l246_6) begin
            if(when_ArraySlice_l276_6) begin
              outputStreamArrayData_6_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l301_6) begin
            outputStreamArrayData_6_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_6_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            outputStreamArrayData_6_payload = _zz_outputStreamArrayData_6_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            outputStreamArrayData_6_payload = _zz_outputStreamArrayData_6_payload_1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_7_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            outputStreamArrayData_7_valid = _zz_outputStreamArrayData_7_valid_2;
          end
          if(when_ArraySlice_l379_7) begin
            if(when_ArraySlice_l409_7) begin
              outputStreamArrayData_7_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l434_7) begin
            outputStreamArrayData_7_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            outputStreamArrayData_7_valid = _zz_outputStreamArrayData_7_valid_3;
          end
          if(when_ArraySlice_l246_7) begin
            if(when_ArraySlice_l276_7) begin
              outputStreamArrayData_7_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l301_7) begin
            outputStreamArrayData_7_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_7_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            outputStreamArrayData_7_payload = _zz_outputStreamArrayData_7_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            outputStreamArrayData_7_payload = _zz_outputStreamArrayData_7_payload_1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_0_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[0]) begin
            fifoGroup_0_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[0]) begin
              fifoGroup_0_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_0_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[0]) begin
            fifoGroup_0_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[0]) begin
              fifoGroup_0_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_0_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_1_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[1]) begin
            fifoGroup_1_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[1]) begin
              fifoGroup_1_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_1_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[1]) begin
            fifoGroup_1_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[1]) begin
              fifoGroup_1_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_1_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_2_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[2]) begin
            fifoGroup_2_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[2]) begin
              fifoGroup_2_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_2_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[2]) begin
            fifoGroup_2_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[2]) begin
              fifoGroup_2_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_2_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_3_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[3]) begin
            fifoGroup_3_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[3]) begin
              fifoGroup_3_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_3_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[3]) begin
            fifoGroup_3_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[3]) begin
              fifoGroup_3_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_3_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_4_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[4]) begin
            fifoGroup_4_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[4]) begin
              fifoGroup_4_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_4_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[4]) begin
            fifoGroup_4_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[4]) begin
              fifoGroup_4_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_4_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_5_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[5]) begin
            fifoGroup_5_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[5]) begin
              fifoGroup_5_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_5_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[5]) begin
            fifoGroup_5_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[5]) begin
              fifoGroup_5_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_5_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_6_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[6]) begin
            fifoGroup_6_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[6]) begin
              fifoGroup_6_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_6_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[6]) begin
            fifoGroup_6_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[6]) begin
              fifoGroup_6_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_6_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_7_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[7]) begin
            fifoGroup_7_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[7]) begin
              fifoGroup_7_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_7_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[7]) begin
            fifoGroup_7_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[7]) begin
              fifoGroup_7_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_7_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_8_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[8]) begin
            fifoGroup_8_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[8]) begin
              fifoGroup_8_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_8_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[8]) begin
            fifoGroup_8_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[8]) begin
              fifoGroup_8_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_8_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_9_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[9]) begin
            fifoGroup_9_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[9]) begin
              fifoGroup_9_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_9_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[9]) begin
            fifoGroup_9_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[9]) begin
              fifoGroup_9_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_9_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_10_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[10]) begin
            fifoGroup_10_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[10]) begin
              fifoGroup_10_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_10_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[10]) begin
            fifoGroup_10_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[10]) begin
              fifoGroup_10_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_10_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_11_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[11]) begin
            fifoGroup_11_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[11]) begin
              fifoGroup_11_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_11_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[11]) begin
            fifoGroup_11_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[11]) begin
              fifoGroup_11_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_11_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_12_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[12]) begin
            fifoGroup_12_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[12]) begin
              fifoGroup_12_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_12_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[12]) begin
            fifoGroup_12_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[12]) begin
              fifoGroup_12_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_12_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_13_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[13]) begin
            fifoGroup_13_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[13]) begin
              fifoGroup_13_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_13_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[13]) begin
            fifoGroup_13_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[13]) begin
              fifoGroup_13_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_13_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_14_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[14]) begin
            fifoGroup_14_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[14]) begin
              fifoGroup_14_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_14_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[14]) begin
            fifoGroup_14_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[14]) begin
              fifoGroup_14_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_14_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_15_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[15]) begin
            fifoGroup_15_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[15]) begin
              fifoGroup_15_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_15_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[15]) begin
            fifoGroup_15_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[15]) begin
              fifoGroup_15_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_15_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_16_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[16]) begin
            fifoGroup_16_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[16]) begin
              fifoGroup_16_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_16_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[16]) begin
            fifoGroup_16_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[16]) begin
              fifoGroup_16_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_16_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_17_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[17]) begin
            fifoGroup_17_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[17]) begin
              fifoGroup_17_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_17_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[17]) begin
            fifoGroup_17_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[17]) begin
              fifoGroup_17_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_17_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_18_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[18]) begin
            fifoGroup_18_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[18]) begin
              fifoGroup_18_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_18_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[18]) begin
            fifoGroup_18_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[18]) begin
              fifoGroup_18_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_18_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_19_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[19]) begin
            fifoGroup_19_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[19]) begin
              fifoGroup_19_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_19_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[19]) begin
            fifoGroup_19_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[19]) begin
              fifoGroup_19_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_19_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_20_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[20]) begin
            fifoGroup_20_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[20]) begin
              fifoGroup_20_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_20_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[20]) begin
            fifoGroup_20_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[20]) begin
              fifoGroup_20_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_20_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_21_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[21]) begin
            fifoGroup_21_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[21]) begin
              fifoGroup_21_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_21_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[21]) begin
            fifoGroup_21_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[21]) begin
              fifoGroup_21_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_21_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_22_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[22]) begin
            fifoGroup_22_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[22]) begin
              fifoGroup_22_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_22_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[22]) begin
            fifoGroup_22_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[22]) begin
              fifoGroup_22_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_22_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_23_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[23]) begin
            fifoGroup_23_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[23]) begin
              fifoGroup_23_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_23_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[23]) begin
            fifoGroup_23_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[23]) begin
              fifoGroup_23_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_23_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_24_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[24]) begin
            fifoGroup_24_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[24]) begin
              fifoGroup_24_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_24_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[24]) begin
            fifoGroup_24_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[24]) begin
              fifoGroup_24_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_24_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_25_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[25]) begin
            fifoGroup_25_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[25]) begin
              fifoGroup_25_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_25_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[25]) begin
            fifoGroup_25_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[25]) begin
              fifoGroup_25_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_25_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_26_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[26]) begin
            fifoGroup_26_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[26]) begin
              fifoGroup_26_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_26_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[26]) begin
            fifoGroup_26_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[26]) begin
              fifoGroup_26_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_26_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_27_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[27]) begin
            fifoGroup_27_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[27]) begin
              fifoGroup_27_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_27_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[27]) begin
            fifoGroup_27_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[27]) begin
              fifoGroup_27_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_27_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_28_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[28]) begin
            fifoGroup_28_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[28]) begin
              fifoGroup_28_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_28_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[28]) begin
            fifoGroup_28_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[28]) begin
              fifoGroup_28_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_28_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_29_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[29]) begin
            fifoGroup_29_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[29]) begin
              fifoGroup_29_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_29_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[29]) begin
            fifoGroup_29_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[29]) begin
              fifoGroup_29_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_29_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_30_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[30]) begin
            fifoGroup_30_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[30]) begin
              fifoGroup_30_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_30_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[30]) begin
            fifoGroup_30_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[30]) begin
              fifoGroup_30_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_30_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_31_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[31]) begin
            fifoGroup_31_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[31]) begin
              fifoGroup_31_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_31_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[31]) begin
            fifoGroup_31_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[31]) begin
              fifoGroup_31_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_31_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_32_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[32]) begin
            fifoGroup_32_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[32]) begin
              fifoGroup_32_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_32_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[32]) begin
            fifoGroup_32_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[32]) begin
              fifoGroup_32_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_32_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_33_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[33]) begin
            fifoGroup_33_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[33]) begin
              fifoGroup_33_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_33_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[33]) begin
            fifoGroup_33_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[33]) begin
              fifoGroup_33_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_33_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_34_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[34]) begin
            fifoGroup_34_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[34]) begin
              fifoGroup_34_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_34_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[34]) begin
            fifoGroup_34_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[34]) begin
              fifoGroup_34_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_34_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_35_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[35]) begin
            fifoGroup_35_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[35]) begin
              fifoGroup_35_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_35_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[35]) begin
            fifoGroup_35_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[35]) begin
              fifoGroup_35_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_35_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_36_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[36]) begin
            fifoGroup_36_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[36]) begin
              fifoGroup_36_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_36_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[36]) begin
            fifoGroup_36_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[36]) begin
              fifoGroup_36_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_36_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_37_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[37]) begin
            fifoGroup_37_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[37]) begin
              fifoGroup_37_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_37_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[37]) begin
            fifoGroup_37_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[37]) begin
              fifoGroup_37_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_37_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_38_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[38]) begin
            fifoGroup_38_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[38]) begin
              fifoGroup_38_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_38_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[38]) begin
            fifoGroup_38_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[38]) begin
              fifoGroup_38_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_38_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_39_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[39]) begin
            fifoGroup_39_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[39]) begin
              fifoGroup_39_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_39_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[39]) begin
            fifoGroup_39_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[39]) begin
              fifoGroup_39_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_39_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_40_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[40]) begin
            fifoGroup_40_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[40]) begin
              fifoGroup_40_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_40_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[40]) begin
            fifoGroup_40_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[40]) begin
              fifoGroup_40_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_40_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_41_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[41]) begin
            fifoGroup_41_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[41]) begin
              fifoGroup_41_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_41_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[41]) begin
            fifoGroup_41_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[41]) begin
              fifoGroup_41_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_41_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_42_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[42]) begin
            fifoGroup_42_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[42]) begin
              fifoGroup_42_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_42_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[42]) begin
            fifoGroup_42_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[42]) begin
              fifoGroup_42_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_42_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_43_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[43]) begin
            fifoGroup_43_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[43]) begin
              fifoGroup_43_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_43_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[43]) begin
            fifoGroup_43_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[43]) begin
              fifoGroup_43_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_43_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_44_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[44]) begin
            fifoGroup_44_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[44]) begin
              fifoGroup_44_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_44_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[44]) begin
            fifoGroup_44_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[44]) begin
              fifoGroup_44_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_44_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_45_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[45]) begin
            fifoGroup_45_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[45]) begin
              fifoGroup_45_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_45_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[45]) begin
            fifoGroup_45_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[45]) begin
              fifoGroup_45_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_45_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_46_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[46]) begin
            fifoGroup_46_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[46]) begin
              fifoGroup_46_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_46_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[46]) begin
            fifoGroup_46_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[46]) begin
              fifoGroup_46_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_46_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_47_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[47]) begin
            fifoGroup_47_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[47]) begin
              fifoGroup_47_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_47_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[47]) begin
            fifoGroup_47_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[47]) begin
              fifoGroup_47_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_47_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_48_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[48]) begin
            fifoGroup_48_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[48]) begin
              fifoGroup_48_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_48_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[48]) begin
            fifoGroup_48_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[48]) begin
              fifoGroup_48_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_48_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_49_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[49]) begin
            fifoGroup_49_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[49]) begin
              fifoGroup_49_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_49_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[49]) begin
            fifoGroup_49_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[49]) begin
              fifoGroup_49_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_49_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_50_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[50]) begin
            fifoGroup_50_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[50]) begin
              fifoGroup_50_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_50_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[50]) begin
            fifoGroup_50_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[50]) begin
              fifoGroup_50_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_50_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_51_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[51]) begin
            fifoGroup_51_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[51]) begin
              fifoGroup_51_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_51_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[51]) begin
            fifoGroup_51_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[51]) begin
              fifoGroup_51_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_51_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_52_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[52]) begin
            fifoGroup_52_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[52]) begin
              fifoGroup_52_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_52_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[52]) begin
            fifoGroup_52_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[52]) begin
              fifoGroup_52_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_52_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_53_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[53]) begin
            fifoGroup_53_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[53]) begin
              fifoGroup_53_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_53_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[53]) begin
            fifoGroup_53_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[53]) begin
              fifoGroup_53_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_53_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_54_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[54]) begin
            fifoGroup_54_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[54]) begin
              fifoGroup_54_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_54_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[54]) begin
            fifoGroup_54_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[54]) begin
              fifoGroup_54_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_54_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_55_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[55]) begin
            fifoGroup_55_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[55]) begin
              fifoGroup_55_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_55_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[55]) begin
            fifoGroup_55_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[55]) begin
              fifoGroup_55_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_55_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_56_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[56]) begin
            fifoGroup_56_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[56]) begin
              fifoGroup_56_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_56_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[56]) begin
            fifoGroup_56_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[56]) begin
              fifoGroup_56_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_56_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_57_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[57]) begin
            fifoGroup_57_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[57]) begin
              fifoGroup_57_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_57_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[57]) begin
            fifoGroup_57_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[57]) begin
              fifoGroup_57_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_57_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_58_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[58]) begin
            fifoGroup_58_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[58]) begin
              fifoGroup_58_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_58_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[58]) begin
            fifoGroup_58_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[58]) begin
              fifoGroup_58_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_58_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_59_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[59]) begin
            fifoGroup_59_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[59]) begin
              fifoGroup_59_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_59_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[59]) begin
            fifoGroup_59_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[59]) begin
              fifoGroup_59_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_59_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_60_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[60]) begin
            fifoGroup_60_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[60]) begin
              fifoGroup_60_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_60_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[60]) begin
            fifoGroup_60_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[60]) begin
              fifoGroup_60_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_60_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_61_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[61]) begin
            fifoGroup_61_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[61]) begin
              fifoGroup_61_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_61_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[61]) begin
            fifoGroup_61_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[61]) begin
              fifoGroup_61_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_61_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_62_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[62]) begin
            fifoGroup_62_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[62]) begin
              fifoGroup_62_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_62_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[62]) begin
            fifoGroup_62_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[62]) begin
              fifoGroup_62_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_62_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_63_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_1[63]) begin
            fifoGroup_63_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_19[63]) begin
              fifoGroup_63_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_63_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l211) begin
          if(_zz_2[63]) begin
            fifoGroup_63_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l333) begin
          if(when_ArraySlice_l334) begin
            if(_zz_20[63]) begin
              fifoGroup_63_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_63_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l373) begin
          if(when_ArraySlice_l374) begin
            if(_zz_3[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l373_1) begin
          if(when_ArraySlice_l374_1) begin
            if(_zz_4[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l373_2) begin
          if(when_ArraySlice_l374_2) begin
            if(_zz_5[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l373_3) begin
          if(when_ArraySlice_l374_3) begin
            if(_zz_6[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l373_4) begin
          if(when_ArraySlice_l374_4) begin
            if(_zz_7[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l373_5) begin
          if(when_ArraySlice_l374_5) begin
            if(_zz_8[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l373_6) begin
          if(when_ArraySlice_l374_6) begin
            if(_zz_9[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l373_7) begin
          if(when_ArraySlice_l374_7) begin
            if(_zz_10[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l240) begin
          if(when_ArraySlice_l241) begin
            if(_zz_11[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l240_1) begin
          if(when_ArraySlice_l241_1) begin
            if(_zz_12[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l240_2) begin
          if(when_ArraySlice_l241_2) begin
            if(_zz_13[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l240_3) begin
          if(when_ArraySlice_l241_3) begin
            if(_zz_14[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l240_4) begin
          if(when_ArraySlice_l241_4) begin
            if(_zz_15[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l240_5) begin
          if(when_ArraySlice_l241_5) begin
            if(_zz_16[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l240_6) begin
          if(when_ArraySlice_l241_6) begin
            if(_zz_17[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l240_7) begin
          if(when_ArraySlice_l241_7) begin
            if(_zz_18[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign arraySliceStateMachine_wantExit = 1'b0;
  always @(*) begin
    arraySliceStateMachine_wantStart = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
      end
      default : begin
        arraySliceStateMachine_wantStart = 1'b1;
      end
    endcase
  end

  assign arraySliceStateMachine_wantKill = 1'b0;
  always @(*) begin
    arraySliceStateMachine_stateNext = arraySliceStateMachine_stateReg;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l223) begin
          arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_readWriteData;
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l465) begin
          arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_readWriteData;
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l354) begin
          arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_writeDataOnly;
        end
        if(when_ArraySlice_l358) begin
          arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_readDataOnly;
        end
      end
      default : begin
      end
    endcase
    if(arraySliceStateMachine_wantStart) begin
      arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_writeDataOnly;
    end
    if(arraySliceStateMachine_wantKill) begin
      arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_BOOT;
    end
  end

  assign when_ArraySlice_l211 = (_zz_when_ArraySlice_l211 < _zz_when_ArraySlice_l211_1);
  assign _zz_1 = ({63'd0,1'b1} <<< selectWriteFifo);
  assign _zz_2 = ({63'd0,1'b1} <<< selectWriteFifo);
  assign _zz_io_push_valid = inputStreamArrayData_valid;
  assign _zz_io_push_payload = inputStreamArrayData_payload;
  assign inputStreamArrayData_fire = (inputStreamArrayData_valid && inputStreamArrayData_ready);
  assign when_ArraySlice_l215 = ((_zz_when_ArraySlice_l215 == _zz_when_ArraySlice_l215_1) && inputStreamArrayData_fire);
  assign when_ArraySlice_l216 = (selectWriteFifo == _zz_when_ArraySlice_l216);
  always @(*) begin
    debug_0 = 1'b0;
    if(when_ArraySlice_l165) begin
      if(when_ArraySlice_l166) begin
        debug_0 = 1'b1;
      end else begin
        debug_0 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173) begin
        debug_0 = 1'b1;
      end else begin
        debug_0 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1 = 1'b0;
    if(when_ArraySlice_l165_1) begin
      if(when_ArraySlice_l166_1) begin
        debug_1 = 1'b1;
      end else begin
        debug_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_1) begin
        debug_1 = 1'b1;
      end else begin
        debug_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2 = 1'b0;
    if(when_ArraySlice_l165_2) begin
      if(when_ArraySlice_l166_2) begin
        debug_2 = 1'b1;
      end else begin
        debug_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_2) begin
        debug_2 = 1'b1;
      end else begin
        debug_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3 = 1'b0;
    if(when_ArraySlice_l165_3) begin
      if(when_ArraySlice_l166_3) begin
        debug_3 = 1'b1;
      end else begin
        debug_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_3) begin
        debug_3 = 1'b1;
      end else begin
        debug_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4 = 1'b0;
    if(when_ArraySlice_l165_4) begin
      if(when_ArraySlice_l166_4) begin
        debug_4 = 1'b1;
      end else begin
        debug_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_4) begin
        debug_4 = 1'b1;
      end else begin
        debug_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5 = 1'b0;
    if(when_ArraySlice_l165_5) begin
      if(when_ArraySlice_l166_5) begin
        debug_5 = 1'b1;
      end else begin
        debug_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_5) begin
        debug_5 = 1'b1;
      end else begin
        debug_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6 = 1'b0;
    if(when_ArraySlice_l165_6) begin
      if(when_ArraySlice_l166_6) begin
        debug_6 = 1'b1;
      end else begin
        debug_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_6) begin
        debug_6 = 1'b1;
      end else begin
        debug_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7 = 1'b0;
    if(when_ArraySlice_l165_7) begin
      if(when_ArraySlice_l166_7) begin
        debug_7 = 1'b1;
      end else begin
        debug_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_7) begin
        debug_7 = 1'b1;
      end else begin
        debug_7 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165 = (_zz_when_ArraySlice_l165 <= selectWriteFifo);
  assign when_ArraySlice_l166 = (_zz_when_ArraySlice_l166 <= _zz_when_ArraySlice_l166_1);
  assign _zz_when_ArraySlice_l112 = (wReg % _zz__zz_when_ArraySlice_l112);
  assign when_ArraySlice_l112 = (_zz_when_ArraySlice_l112 != 6'h0);
  assign when_ArraySlice_l113 = (7'h40 <= _zz_when_ArraySlice_l113);
  always @(*) begin
    if(when_ArraySlice_l112) begin
      if(when_ArraySlice_l113) begin
        _zz_when_ArraySlice_l173 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173 = (_zz__zz_when_ArraySlice_l173 - _zz__zz_when_ArraySlice_l173_3);
      end
    end else begin
      if(when_ArraySlice_l118) begin
        _zz_when_ArraySlice_l173 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118 = (_zz_when_ArraySlice_l118 <= wReg);
  assign when_ArraySlice_l173 = (_zz_when_ArraySlice_l173_416 <= _zz_when_ArraySlice_l173_417);
  assign when_ArraySlice_l165_1 = (_zz_when_ArraySlice_l165_1_1 <= selectWriteFifo);
  assign when_ArraySlice_l166_1 = (_zz_when_ArraySlice_l166_1_1 <= _zz_when_ArraySlice_l166_1_2);
  assign _zz_when_ArraySlice_l112_1 = (wReg % _zz__zz_when_ArraySlice_l112_1);
  assign when_ArraySlice_l112_1 = (_zz_when_ArraySlice_l112_1 != 6'h0);
  assign when_ArraySlice_l113_1 = (7'h40 <= _zz_when_ArraySlice_l113_1_1);
  always @(*) begin
    if(when_ArraySlice_l112_1) begin
      if(when_ArraySlice_l113_1) begin
        _zz_when_ArraySlice_l173_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_1 = (_zz__zz_when_ArraySlice_l173_1_1 - _zz__zz_when_ArraySlice_l173_1_4);
      end
    end else begin
      if(when_ArraySlice_l118_1) begin
        _zz_when_ArraySlice_l173_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_1 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_1 = (_zz_when_ArraySlice_l118_1_1 <= wReg);
  assign when_ArraySlice_l173_1 = (_zz_when_ArraySlice_l173_1_1 <= _zz_when_ArraySlice_l173_1_3);
  assign when_ArraySlice_l165_2 = (_zz_when_ArraySlice_l165_2_1 <= selectWriteFifo);
  assign when_ArraySlice_l166_2 = (_zz_when_ArraySlice_l166_2_1 <= _zz_when_ArraySlice_l166_2_2);
  assign _zz_when_ArraySlice_l112_2 = (wReg % _zz__zz_when_ArraySlice_l112_2);
  assign when_ArraySlice_l112_2 = (_zz_when_ArraySlice_l112_2 != 6'h0);
  assign when_ArraySlice_l113_2 = (7'h40 <= _zz_when_ArraySlice_l113_2_1);
  always @(*) begin
    if(when_ArraySlice_l112_2) begin
      if(when_ArraySlice_l113_2) begin
        _zz_when_ArraySlice_l173_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_2 = (_zz__zz_when_ArraySlice_l173_2_1 - _zz__zz_when_ArraySlice_l173_2_4);
      end
    end else begin
      if(when_ArraySlice_l118_2) begin
        _zz_when_ArraySlice_l173_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_2 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_2 = (_zz_when_ArraySlice_l118_2 <= wReg);
  assign when_ArraySlice_l173_2 = (_zz_when_ArraySlice_l173_2_1 <= _zz_when_ArraySlice_l173_2_3);
  assign when_ArraySlice_l165_3 = (_zz_when_ArraySlice_l165_3 <= selectWriteFifo);
  assign when_ArraySlice_l166_3 = (_zz_when_ArraySlice_l166_3_1 <= _zz_when_ArraySlice_l166_3_2);
  assign _zz_when_ArraySlice_l112_3 = (wReg % _zz__zz_when_ArraySlice_l112_3);
  assign when_ArraySlice_l112_3 = (_zz_when_ArraySlice_l112_3 != 6'h0);
  assign when_ArraySlice_l113_3 = (7'h40 <= _zz_when_ArraySlice_l113_3_1);
  always @(*) begin
    if(when_ArraySlice_l112_3) begin
      if(when_ArraySlice_l113_3) begin
        _zz_when_ArraySlice_l173_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_3 = (_zz__zz_when_ArraySlice_l173_3_1 - _zz__zz_when_ArraySlice_l173_3_4);
      end
    end else begin
      if(when_ArraySlice_l118_3) begin
        _zz_when_ArraySlice_l173_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_3 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_3 = (_zz_when_ArraySlice_l118_3 <= wReg);
  assign when_ArraySlice_l173_3 = (_zz_when_ArraySlice_l173_3_1 <= _zz_when_ArraySlice_l173_3_3);
  assign when_ArraySlice_l165_4 = (_zz_when_ArraySlice_l165_4 <= selectWriteFifo);
  assign when_ArraySlice_l166_4 = (_zz_when_ArraySlice_l166_4_1 <= _zz_when_ArraySlice_l166_4_2);
  assign _zz_when_ArraySlice_l112_4 = (wReg % _zz__zz_when_ArraySlice_l112_4);
  assign when_ArraySlice_l112_4 = (_zz_when_ArraySlice_l112_4 != 6'h0);
  assign when_ArraySlice_l113_4 = (7'h40 <= _zz_when_ArraySlice_l113_4_1);
  always @(*) begin
    if(when_ArraySlice_l112_4) begin
      if(when_ArraySlice_l113_4) begin
        _zz_when_ArraySlice_l173_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_4 = (_zz__zz_when_ArraySlice_l173_4 - _zz__zz_when_ArraySlice_l173_4_3);
      end
    end else begin
      if(when_ArraySlice_l118_4) begin
        _zz_when_ArraySlice_l173_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_4 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_4 = (_zz_when_ArraySlice_l118_4 <= wReg);
  assign when_ArraySlice_l173_4 = (_zz_when_ArraySlice_l173_4_1 <= _zz_when_ArraySlice_l173_4_3);
  assign when_ArraySlice_l165_5 = (_zz_when_ArraySlice_l165_5 <= selectWriteFifo);
  assign when_ArraySlice_l166_5 = (_zz_when_ArraySlice_l166_5_1 <= _zz_when_ArraySlice_l166_5_3);
  assign _zz_when_ArraySlice_l112_5 = (wReg % _zz__zz_when_ArraySlice_l112_5);
  assign when_ArraySlice_l112_5 = (_zz_when_ArraySlice_l112_5 != 6'h0);
  assign when_ArraySlice_l113_5 = (7'h40 <= _zz_when_ArraySlice_l113_5);
  always @(*) begin
    if(when_ArraySlice_l112_5) begin
      if(when_ArraySlice_l113_5) begin
        _zz_when_ArraySlice_l173_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_5 = (_zz__zz_when_ArraySlice_l173_5 - _zz__zz_when_ArraySlice_l173_5_3);
      end
    end else begin
      if(when_ArraySlice_l118_5) begin
        _zz_when_ArraySlice_l173_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_5 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_5 = (_zz_when_ArraySlice_l118_5 <= wReg);
  assign when_ArraySlice_l173_5 = (_zz_when_ArraySlice_l173_5_1 <= _zz_when_ArraySlice_l173_5_3);
  assign when_ArraySlice_l165_6 = (_zz_when_ArraySlice_l165_6 <= selectWriteFifo);
  assign when_ArraySlice_l166_6 = (_zz_when_ArraySlice_l166_6 <= _zz_when_ArraySlice_l166_6_2);
  assign _zz_when_ArraySlice_l112_6 = (wReg % _zz__zz_when_ArraySlice_l112_6);
  assign when_ArraySlice_l112_6 = (_zz_when_ArraySlice_l112_6 != 6'h0);
  assign when_ArraySlice_l113_6 = (7'h40 <= _zz_when_ArraySlice_l113_6);
  always @(*) begin
    if(when_ArraySlice_l112_6) begin
      if(when_ArraySlice_l113_6) begin
        _zz_when_ArraySlice_l173_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_6 = (_zz__zz_when_ArraySlice_l173_6 - _zz__zz_when_ArraySlice_l173_6_3);
      end
    end else begin
      if(when_ArraySlice_l118_6) begin
        _zz_when_ArraySlice_l173_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_6 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_6 = (_zz_when_ArraySlice_l118_6 <= wReg);
  assign when_ArraySlice_l173_6 = (_zz_when_ArraySlice_l173_6_1 <= _zz_when_ArraySlice_l173_6_3);
  assign when_ArraySlice_l165_7 = (_zz_when_ArraySlice_l165_7 <= selectWriteFifo);
  assign when_ArraySlice_l166_7 = (_zz_when_ArraySlice_l166_7 <= _zz_when_ArraySlice_l166_7_2);
  assign _zz_when_ArraySlice_l112_7 = (wReg % _zz__zz_when_ArraySlice_l112_7);
  assign when_ArraySlice_l112_7 = (_zz_when_ArraySlice_l112_7 != 6'h0);
  assign when_ArraySlice_l113_7 = (7'h40 <= _zz_when_ArraySlice_l113_7);
  always @(*) begin
    if(when_ArraySlice_l112_7) begin
      if(when_ArraySlice_l113_7) begin
        _zz_when_ArraySlice_l173_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_7 = (_zz__zz_when_ArraySlice_l173_7 - _zz__zz_when_ArraySlice_l173_7_3);
      end
    end else begin
      if(when_ArraySlice_l118_7) begin
        _zz_when_ArraySlice_l173_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_7 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_7 = (_zz_when_ArraySlice_l118_7 <= wReg);
  assign when_ArraySlice_l173_7 = (_zz_when_ArraySlice_l173_7_1 <= _zz_when_ArraySlice_l173_7_3);
  assign when_ArraySlice_l223 = ((((((((debug_0 == 1'b1) && (debug_1 == 1'b1)) && (debug_2 == 1'b1)) && (debug_3 == 1'b1)) && (debug_4 == 1'b1)) && (debug_5 == 1'b1)) && (debug_6 == 1'b1)) && (debug_7 == 1'b1));
  assign when_ArraySlice_l229 = (! allowPadding_0);
  assign when_ArraySlice_l229_1 = (! allowPadding_1);
  assign when_ArraySlice_l229_2 = (! allowPadding_2);
  assign when_ArraySlice_l229_3 = (! allowPadding_3);
  assign when_ArraySlice_l229_4 = (! allowPadding_4);
  assign when_ArraySlice_l229_5 = (! allowPadding_5);
  assign when_ArraySlice_l229_6 = (! allowPadding_6);
  assign when_ArraySlice_l229_7 = (! allowPadding_7);
  assign when_ArraySlice_l373 = (_zz_when_ArraySlice_l373 < wReg);
  assign when_ArraySlice_l374 = ((! holdReadOp_0) && (_zz_when_ArraySlice_l374 != 7'h0));
  assign _zz_outputStreamArrayData_0_valid = (selectReadFifo_0 + _zz__zz_outputStreamArrayData_0_valid);
  assign _zz_3 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_0_valid);
  assign _zz_io_pop_ready = outputStreamArrayData_0_ready;
  assign when_ArraySlice_l379 = (! holdReadOp_0);
  assign outputStreamArrayData_0_fire = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l380 = ((_zz_when_ArraySlice_l380 < _zz_when_ArraySlice_l380_2) && outputStreamArrayData_0_fire);
  assign when_ArraySlice_l381 = (handshakeTimes_0_value == _zz_when_ArraySlice_l381);
  assign when_ArraySlice_l384 = (_zz_when_ArraySlice_l384 == 13'h0);
  assign outputStreamArrayData_0_fire_1 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l389 = ((_zz_when_ArraySlice_l389 == _zz_when_ArraySlice_l389_4) && outputStreamArrayData_0_fire_1);
  assign when_ArraySlice_l390 = (handshakeTimes_0_value == _zz_when_ArraySlice_l390);
  assign _zz_when_ArraySlice_l94 = (hReg % _zz__zz_when_ArraySlice_l94);
  assign when_ArraySlice_l94 = (_zz_when_ArraySlice_l94 != 6'h0);
  assign when_ArraySlice_l95 = (7'h40 <= _zz_when_ArraySlice_l95);
  always @(*) begin
    if(when_ArraySlice_l94) begin
      if(when_ArraySlice_l95) begin
        _zz_when_ArraySlice_l392 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392 = (_zz__zz_when_ArraySlice_l392 - _zz__zz_when_ArraySlice_l392_3);
      end
    end else begin
      if(when_ArraySlice_l99) begin
        _zz_when_ArraySlice_l392 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99 = (_zz_when_ArraySlice_l99 <= hReg);
  assign when_ArraySlice_l392 = (_zz_when_ArraySlice_l392_8 < _zz_when_ArraySlice_l392_11);
  always @(*) begin
    debug_0_1 = 1'b0;
    if(when_ArraySlice_l165_8) begin
      if(when_ArraySlice_l166_8) begin
        debug_0_1 = 1'b1;
      end else begin
        debug_0_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_8) begin
        debug_0_1 = 1'b1;
      end else begin
        debug_0_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_1 = 1'b0;
    if(when_ArraySlice_l165_9) begin
      if(when_ArraySlice_l166_9) begin
        debug_1_1 = 1'b1;
      end else begin
        debug_1_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_9) begin
        debug_1_1 = 1'b1;
      end else begin
        debug_1_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_1 = 1'b0;
    if(when_ArraySlice_l165_10) begin
      if(when_ArraySlice_l166_10) begin
        debug_2_1 = 1'b1;
      end else begin
        debug_2_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_10) begin
        debug_2_1 = 1'b1;
      end else begin
        debug_2_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_1 = 1'b0;
    if(when_ArraySlice_l165_11) begin
      if(when_ArraySlice_l166_11) begin
        debug_3_1 = 1'b1;
      end else begin
        debug_3_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_11) begin
        debug_3_1 = 1'b1;
      end else begin
        debug_3_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_1 = 1'b0;
    if(when_ArraySlice_l165_12) begin
      if(when_ArraySlice_l166_12) begin
        debug_4_1 = 1'b1;
      end else begin
        debug_4_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_12) begin
        debug_4_1 = 1'b1;
      end else begin
        debug_4_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_1 = 1'b0;
    if(when_ArraySlice_l165_13) begin
      if(when_ArraySlice_l166_13) begin
        debug_5_1 = 1'b1;
      end else begin
        debug_5_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_13) begin
        debug_5_1 = 1'b1;
      end else begin
        debug_5_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_1 = 1'b0;
    if(when_ArraySlice_l165_14) begin
      if(when_ArraySlice_l166_14) begin
        debug_6_1 = 1'b1;
      end else begin
        debug_6_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_14) begin
        debug_6_1 = 1'b1;
      end else begin
        debug_6_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_1 = 1'b0;
    if(when_ArraySlice_l165_15) begin
      if(when_ArraySlice_l166_15) begin
        debug_7_1 = 1'b1;
      end else begin
        debug_7_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_15) begin
        debug_7_1 = 1'b1;
      end else begin
        debug_7_1 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_8 = (_zz_when_ArraySlice_l165_8 <= selectWriteFifo);
  assign when_ArraySlice_l166_8 = (_zz_when_ArraySlice_l166_8 <= _zz_when_ArraySlice_l166_8_1);
  assign _zz_when_ArraySlice_l112_8 = (wReg % _zz__zz_when_ArraySlice_l112_8);
  assign when_ArraySlice_l112_8 = (_zz_when_ArraySlice_l112_8 != 6'h0);
  assign when_ArraySlice_l113_8 = (7'h40 <= _zz_when_ArraySlice_l113_8);
  always @(*) begin
    if(when_ArraySlice_l112_8) begin
      if(when_ArraySlice_l113_8) begin
        _zz_when_ArraySlice_l173_8 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_8 = (_zz__zz_when_ArraySlice_l173_8 - _zz__zz_when_ArraySlice_l173_8_3);
      end
    end else begin
      if(when_ArraySlice_l118_8) begin
        _zz_when_ArraySlice_l173_8 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_8 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_8 = (_zz_when_ArraySlice_l118_8 <= wReg);
  assign when_ArraySlice_l173_8 = (_zz_when_ArraySlice_l173_8_1 <= _zz_when_ArraySlice_l173_8_2);
  assign when_ArraySlice_l165_9 = (_zz_when_ArraySlice_l165_9 <= selectWriteFifo);
  assign when_ArraySlice_l166_9 = (_zz_when_ArraySlice_l166_9 <= _zz_when_ArraySlice_l166_9_1);
  assign _zz_when_ArraySlice_l112_9 = (wReg % _zz__zz_when_ArraySlice_l112_9);
  assign when_ArraySlice_l112_9 = (_zz_when_ArraySlice_l112_9 != 6'h0);
  assign when_ArraySlice_l113_9 = (7'h40 <= _zz_when_ArraySlice_l113_9);
  always @(*) begin
    if(when_ArraySlice_l112_9) begin
      if(when_ArraySlice_l113_9) begin
        _zz_when_ArraySlice_l173_9 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_9 = (_zz__zz_when_ArraySlice_l173_9 - _zz__zz_when_ArraySlice_l173_9_3);
      end
    end else begin
      if(when_ArraySlice_l118_9) begin
        _zz_when_ArraySlice_l173_9 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_9 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_9 = (_zz_when_ArraySlice_l118_9 <= wReg);
  assign when_ArraySlice_l173_9 = (_zz_when_ArraySlice_l173_9_1 <= _zz_when_ArraySlice_l173_9_3);
  assign when_ArraySlice_l165_10 = (_zz_when_ArraySlice_l165_10 <= selectWriteFifo);
  assign when_ArraySlice_l166_10 = (_zz_when_ArraySlice_l166_10 <= _zz_when_ArraySlice_l166_10_1);
  assign _zz_when_ArraySlice_l112_10 = (wReg % _zz__zz_when_ArraySlice_l112_10);
  assign when_ArraySlice_l112_10 = (_zz_when_ArraySlice_l112_10 != 6'h0);
  assign when_ArraySlice_l113_10 = (7'h40 <= _zz_when_ArraySlice_l113_10);
  always @(*) begin
    if(when_ArraySlice_l112_10) begin
      if(when_ArraySlice_l113_10) begin
        _zz_when_ArraySlice_l173_10 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_10 = (_zz__zz_when_ArraySlice_l173_10 - _zz__zz_when_ArraySlice_l173_10_3);
      end
    end else begin
      if(when_ArraySlice_l118_10) begin
        _zz_when_ArraySlice_l173_10 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_10 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_10 = (_zz_when_ArraySlice_l118_10 <= wReg);
  assign when_ArraySlice_l173_10 = (_zz_when_ArraySlice_l173_10_1 <= _zz_when_ArraySlice_l173_10_3);
  assign when_ArraySlice_l165_11 = (_zz_when_ArraySlice_l165_11 <= selectWriteFifo);
  assign when_ArraySlice_l166_11 = (_zz_when_ArraySlice_l166_11 <= _zz_when_ArraySlice_l166_11_1);
  assign _zz_when_ArraySlice_l112_11 = (wReg % _zz__zz_when_ArraySlice_l112_11);
  assign when_ArraySlice_l112_11 = (_zz_when_ArraySlice_l112_11 != 6'h0);
  assign when_ArraySlice_l113_11 = (7'h40 <= _zz_when_ArraySlice_l113_11);
  always @(*) begin
    if(when_ArraySlice_l112_11) begin
      if(when_ArraySlice_l113_11) begin
        _zz_when_ArraySlice_l173_11 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_11 = (_zz__zz_when_ArraySlice_l173_11 - _zz__zz_when_ArraySlice_l173_11_3);
      end
    end else begin
      if(when_ArraySlice_l118_11) begin
        _zz_when_ArraySlice_l173_11 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_11 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_11 = (_zz_when_ArraySlice_l118_11 <= wReg);
  assign when_ArraySlice_l173_11 = (_zz_when_ArraySlice_l173_11_1 <= _zz_when_ArraySlice_l173_11_3);
  assign when_ArraySlice_l165_12 = (_zz_when_ArraySlice_l165_12 <= selectWriteFifo);
  assign when_ArraySlice_l166_12 = (_zz_when_ArraySlice_l166_12 <= _zz_when_ArraySlice_l166_12_1);
  assign _zz_when_ArraySlice_l112_12 = (wReg % _zz__zz_when_ArraySlice_l112_12);
  assign when_ArraySlice_l112_12 = (_zz_when_ArraySlice_l112_12 != 6'h0);
  assign when_ArraySlice_l113_12 = (7'h40 <= _zz_when_ArraySlice_l113_12);
  always @(*) begin
    if(when_ArraySlice_l112_12) begin
      if(when_ArraySlice_l113_12) begin
        _zz_when_ArraySlice_l173_12 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_12 = (_zz__zz_when_ArraySlice_l173_12 - _zz__zz_when_ArraySlice_l173_12_3);
      end
    end else begin
      if(when_ArraySlice_l118_12) begin
        _zz_when_ArraySlice_l173_12 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_12 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_12 = (_zz_when_ArraySlice_l118_12 <= wReg);
  assign when_ArraySlice_l173_12 = (_zz_when_ArraySlice_l173_12_1 <= _zz_when_ArraySlice_l173_12_3);
  assign when_ArraySlice_l165_13 = (_zz_when_ArraySlice_l165_13 <= selectWriteFifo);
  assign when_ArraySlice_l166_13 = (_zz_when_ArraySlice_l166_13 <= _zz_when_ArraySlice_l166_13_2);
  assign _zz_when_ArraySlice_l112_13 = (wReg % _zz__zz_when_ArraySlice_l112_13);
  assign when_ArraySlice_l112_13 = (_zz_when_ArraySlice_l112_13 != 6'h0);
  assign when_ArraySlice_l113_13 = (7'h40 <= _zz_when_ArraySlice_l113_13);
  always @(*) begin
    if(when_ArraySlice_l112_13) begin
      if(when_ArraySlice_l113_13) begin
        _zz_when_ArraySlice_l173_13 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_13 = (_zz__zz_when_ArraySlice_l173_13 - _zz__zz_when_ArraySlice_l173_13_3);
      end
    end else begin
      if(when_ArraySlice_l118_13) begin
        _zz_when_ArraySlice_l173_13 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_13 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_13 = (_zz_when_ArraySlice_l118_13 <= wReg);
  assign when_ArraySlice_l173_13 = (_zz_when_ArraySlice_l173_13_1 <= _zz_when_ArraySlice_l173_13_3);
  assign when_ArraySlice_l165_14 = (_zz_when_ArraySlice_l165_14 <= selectWriteFifo);
  assign when_ArraySlice_l166_14 = (_zz_when_ArraySlice_l166_14 <= _zz_when_ArraySlice_l166_14_2);
  assign _zz_when_ArraySlice_l112_14 = (wReg % _zz__zz_when_ArraySlice_l112_14);
  assign when_ArraySlice_l112_14 = (_zz_when_ArraySlice_l112_14 != 6'h0);
  assign when_ArraySlice_l113_14 = (7'h40 <= _zz_when_ArraySlice_l113_14);
  always @(*) begin
    if(when_ArraySlice_l112_14) begin
      if(when_ArraySlice_l113_14) begin
        _zz_when_ArraySlice_l173_14 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_14 = (_zz__zz_when_ArraySlice_l173_14 - _zz__zz_when_ArraySlice_l173_14_3);
      end
    end else begin
      if(when_ArraySlice_l118_14) begin
        _zz_when_ArraySlice_l173_14 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_14 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_14 = (_zz_when_ArraySlice_l118_14 <= wReg);
  assign when_ArraySlice_l173_14 = (_zz_when_ArraySlice_l173_14_1 <= _zz_when_ArraySlice_l173_14_3);
  assign when_ArraySlice_l165_15 = (_zz_when_ArraySlice_l165_15 <= selectWriteFifo);
  assign when_ArraySlice_l166_15 = (_zz_when_ArraySlice_l166_15 <= _zz_when_ArraySlice_l166_15_2);
  assign _zz_when_ArraySlice_l112_15 = (wReg % _zz__zz_when_ArraySlice_l112_15);
  assign when_ArraySlice_l112_15 = (_zz_when_ArraySlice_l112_15 != 6'h0);
  assign when_ArraySlice_l113_15 = (7'h40 <= _zz_when_ArraySlice_l113_15);
  always @(*) begin
    if(when_ArraySlice_l112_15) begin
      if(when_ArraySlice_l113_15) begin
        _zz_when_ArraySlice_l173_15 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_15 = (_zz__zz_when_ArraySlice_l173_15 - _zz__zz_when_ArraySlice_l173_15_3);
      end
    end else begin
      if(when_ArraySlice_l118_15) begin
        _zz_when_ArraySlice_l173_15 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_15 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_15 = (_zz_when_ArraySlice_l118_15 <= wReg);
  assign when_ArraySlice_l173_15 = (_zz_when_ArraySlice_l173_15_1 <= _zz_when_ArraySlice_l173_15_3);
  assign when_ArraySlice_l398 = (! (((((_zz_when_ArraySlice_l398 && _zz_when_ArraySlice_l398_3) && (holdReadOp_5 == _zz_when_ArraySlice_l398_4)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && ((((_zz_when_ArraySlice_l398_5 && _zz_when_ArraySlice_l398_8) && (debug_5_1 == _zz_when_ArraySlice_l398_9)) && (debug_6_1 == 1'b1)) && (debug_7_1 == 1'b1))));
  assign when_ArraySlice_l401 = (wReg <= _zz_when_ArraySlice_l401);
  assign when_ArraySlice_l405 = (_zz_when_ArraySlice_l405 == 13'h0);
  assign when_ArraySlice_l409 = (_zz_when_ArraySlice_l409 == 7'h0);
  assign outputStreamArrayData_0_fire_2 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l410 = ((handshakeTimes_0_value == _zz_when_ArraySlice_l410) && outputStreamArrayData_0_fire_2);
  assign _zz_when_ArraySlice_l94_1 = (hReg % _zz__zz_when_ArraySlice_l94_1);
  assign when_ArraySlice_l94_1 = (_zz_when_ArraySlice_l94_1 != 6'h0);
  assign when_ArraySlice_l95_1 = (7'h40 <= _zz_when_ArraySlice_l95_1_1);
  always @(*) begin
    if(when_ArraySlice_l94_1) begin
      if(when_ArraySlice_l95_1) begin
        _zz_when_ArraySlice_l412 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412 = (_zz__zz_when_ArraySlice_l412 - _zz__zz_when_ArraySlice_l412_3);
      end
    end else begin
      if(when_ArraySlice_l99_1) begin
        _zz_when_ArraySlice_l412 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_1 = (_zz_when_ArraySlice_l99_1_1 <= hReg);
  assign when_ArraySlice_l412 = (_zz_when_ArraySlice_l412_8 < _zz_when_ArraySlice_l412_11);
  always @(*) begin
    debug_0_2 = 1'b0;
    if(when_ArraySlice_l165_16) begin
      if(when_ArraySlice_l166_16) begin
        debug_0_2 = 1'b1;
      end else begin
        debug_0_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_16) begin
        debug_0_2 = 1'b1;
      end else begin
        debug_0_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_2 = 1'b0;
    if(when_ArraySlice_l165_17) begin
      if(when_ArraySlice_l166_17) begin
        debug_1_2 = 1'b1;
      end else begin
        debug_1_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_17) begin
        debug_1_2 = 1'b1;
      end else begin
        debug_1_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_2 = 1'b0;
    if(when_ArraySlice_l165_18) begin
      if(when_ArraySlice_l166_18) begin
        debug_2_2 = 1'b1;
      end else begin
        debug_2_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_18) begin
        debug_2_2 = 1'b1;
      end else begin
        debug_2_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_2 = 1'b0;
    if(when_ArraySlice_l165_19) begin
      if(when_ArraySlice_l166_19) begin
        debug_3_2 = 1'b1;
      end else begin
        debug_3_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_19) begin
        debug_3_2 = 1'b1;
      end else begin
        debug_3_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_2 = 1'b0;
    if(when_ArraySlice_l165_20) begin
      if(when_ArraySlice_l166_20) begin
        debug_4_2 = 1'b1;
      end else begin
        debug_4_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_20) begin
        debug_4_2 = 1'b1;
      end else begin
        debug_4_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_2 = 1'b0;
    if(when_ArraySlice_l165_21) begin
      if(when_ArraySlice_l166_21) begin
        debug_5_2 = 1'b1;
      end else begin
        debug_5_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_21) begin
        debug_5_2 = 1'b1;
      end else begin
        debug_5_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_2 = 1'b0;
    if(when_ArraySlice_l165_22) begin
      if(when_ArraySlice_l166_22) begin
        debug_6_2 = 1'b1;
      end else begin
        debug_6_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_22) begin
        debug_6_2 = 1'b1;
      end else begin
        debug_6_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_2 = 1'b0;
    if(when_ArraySlice_l165_23) begin
      if(when_ArraySlice_l166_23) begin
        debug_7_2 = 1'b1;
      end else begin
        debug_7_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_23) begin
        debug_7_2 = 1'b1;
      end else begin
        debug_7_2 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_16 = (_zz_when_ArraySlice_l165_16 <= selectWriteFifo);
  assign when_ArraySlice_l166_16 = (_zz_when_ArraySlice_l166_16 <= _zz_when_ArraySlice_l166_16_1);
  assign _zz_when_ArraySlice_l112_16 = (wReg % _zz__zz_when_ArraySlice_l112_16);
  assign when_ArraySlice_l112_16 = (_zz_when_ArraySlice_l112_16 != 6'h0);
  assign when_ArraySlice_l113_16 = (7'h40 <= _zz_when_ArraySlice_l113_16);
  always @(*) begin
    if(when_ArraySlice_l112_16) begin
      if(when_ArraySlice_l113_16) begin
        _zz_when_ArraySlice_l173_16 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_16 = (_zz__zz_when_ArraySlice_l173_16 - _zz__zz_when_ArraySlice_l173_16_3);
      end
    end else begin
      if(when_ArraySlice_l118_16) begin
        _zz_when_ArraySlice_l173_16 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_16 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_16 = (_zz_when_ArraySlice_l118_16 <= wReg);
  assign when_ArraySlice_l173_16 = (_zz_when_ArraySlice_l173_16_1 <= _zz_when_ArraySlice_l173_16_2);
  assign when_ArraySlice_l165_17 = (_zz_when_ArraySlice_l165_17 <= selectWriteFifo);
  assign when_ArraySlice_l166_17 = (_zz_when_ArraySlice_l166_17 <= _zz_when_ArraySlice_l166_17_1);
  assign _zz_when_ArraySlice_l112_17 = (wReg % _zz__zz_when_ArraySlice_l112_17);
  assign when_ArraySlice_l112_17 = (_zz_when_ArraySlice_l112_17 != 6'h0);
  assign when_ArraySlice_l113_17 = (7'h40 <= _zz_when_ArraySlice_l113_17);
  always @(*) begin
    if(when_ArraySlice_l112_17) begin
      if(when_ArraySlice_l113_17) begin
        _zz_when_ArraySlice_l173_17 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_17 = (_zz__zz_when_ArraySlice_l173_17 - _zz__zz_when_ArraySlice_l173_17_3);
      end
    end else begin
      if(when_ArraySlice_l118_17) begin
        _zz_when_ArraySlice_l173_17 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_17 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_17 = (_zz_when_ArraySlice_l118_17 <= wReg);
  assign when_ArraySlice_l173_17 = (_zz_when_ArraySlice_l173_17_1 <= _zz_when_ArraySlice_l173_17_3);
  assign when_ArraySlice_l165_18 = (_zz_when_ArraySlice_l165_18 <= selectWriteFifo);
  assign when_ArraySlice_l166_18 = (_zz_when_ArraySlice_l166_18 <= _zz_when_ArraySlice_l166_18_1);
  assign _zz_when_ArraySlice_l112_18 = (wReg % _zz__zz_when_ArraySlice_l112_18);
  assign when_ArraySlice_l112_18 = (_zz_when_ArraySlice_l112_18 != 6'h0);
  assign when_ArraySlice_l113_18 = (7'h40 <= _zz_when_ArraySlice_l113_18);
  always @(*) begin
    if(when_ArraySlice_l112_18) begin
      if(when_ArraySlice_l113_18) begin
        _zz_when_ArraySlice_l173_18 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_18 = (_zz__zz_when_ArraySlice_l173_18 - _zz__zz_when_ArraySlice_l173_18_3);
      end
    end else begin
      if(when_ArraySlice_l118_18) begin
        _zz_when_ArraySlice_l173_18 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_18 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_18 = (_zz_when_ArraySlice_l118_18 <= wReg);
  assign when_ArraySlice_l173_18 = (_zz_when_ArraySlice_l173_18_1 <= _zz_when_ArraySlice_l173_18_3);
  assign when_ArraySlice_l165_19 = (_zz_when_ArraySlice_l165_19 <= selectWriteFifo);
  assign when_ArraySlice_l166_19 = (_zz_when_ArraySlice_l166_19 <= _zz_when_ArraySlice_l166_19_1);
  assign _zz_when_ArraySlice_l112_19 = (wReg % _zz__zz_when_ArraySlice_l112_19);
  assign when_ArraySlice_l112_19 = (_zz_when_ArraySlice_l112_19 != 6'h0);
  assign when_ArraySlice_l113_19 = (7'h40 <= _zz_when_ArraySlice_l113_19);
  always @(*) begin
    if(when_ArraySlice_l112_19) begin
      if(when_ArraySlice_l113_19) begin
        _zz_when_ArraySlice_l173_19 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_19 = (_zz__zz_when_ArraySlice_l173_19 - _zz__zz_when_ArraySlice_l173_19_3);
      end
    end else begin
      if(when_ArraySlice_l118_19) begin
        _zz_when_ArraySlice_l173_19 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_19 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_19 = (_zz_when_ArraySlice_l118_19 <= wReg);
  assign when_ArraySlice_l173_19 = (_zz_when_ArraySlice_l173_19_1 <= _zz_when_ArraySlice_l173_19_3);
  assign when_ArraySlice_l165_20 = (_zz_when_ArraySlice_l165_20 <= selectWriteFifo);
  assign when_ArraySlice_l166_20 = (_zz_when_ArraySlice_l166_20 <= _zz_when_ArraySlice_l166_20_1);
  assign _zz_when_ArraySlice_l112_20 = (wReg % _zz__zz_when_ArraySlice_l112_20);
  assign when_ArraySlice_l112_20 = (_zz_when_ArraySlice_l112_20 != 6'h0);
  assign when_ArraySlice_l113_20 = (7'h40 <= _zz_when_ArraySlice_l113_20);
  always @(*) begin
    if(when_ArraySlice_l112_20) begin
      if(when_ArraySlice_l113_20) begin
        _zz_when_ArraySlice_l173_20 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_20 = (_zz__zz_when_ArraySlice_l173_20 - _zz__zz_when_ArraySlice_l173_20_3);
      end
    end else begin
      if(when_ArraySlice_l118_20) begin
        _zz_when_ArraySlice_l173_20 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_20 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_20 = (_zz_when_ArraySlice_l118_20 <= wReg);
  assign when_ArraySlice_l173_20 = (_zz_when_ArraySlice_l173_20_1 <= _zz_when_ArraySlice_l173_20_3);
  assign when_ArraySlice_l165_21 = (_zz_when_ArraySlice_l165_21 <= selectWriteFifo);
  assign when_ArraySlice_l166_21 = (_zz_when_ArraySlice_l166_21 <= _zz_when_ArraySlice_l166_21_2);
  assign _zz_when_ArraySlice_l112_21 = (wReg % _zz__zz_when_ArraySlice_l112_21);
  assign when_ArraySlice_l112_21 = (_zz_when_ArraySlice_l112_21 != 6'h0);
  assign when_ArraySlice_l113_21 = (7'h40 <= _zz_when_ArraySlice_l113_21);
  always @(*) begin
    if(when_ArraySlice_l112_21) begin
      if(when_ArraySlice_l113_21) begin
        _zz_when_ArraySlice_l173_21 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_21 = (_zz__zz_when_ArraySlice_l173_21 - _zz__zz_when_ArraySlice_l173_21_3);
      end
    end else begin
      if(when_ArraySlice_l118_21) begin
        _zz_when_ArraySlice_l173_21 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_21 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_21 = (_zz_when_ArraySlice_l118_21 <= wReg);
  assign when_ArraySlice_l173_21 = (_zz_when_ArraySlice_l173_21_1 <= _zz_when_ArraySlice_l173_21_3);
  assign when_ArraySlice_l165_22 = (_zz_when_ArraySlice_l165_22 <= selectWriteFifo);
  assign when_ArraySlice_l166_22 = (_zz_when_ArraySlice_l166_22 <= _zz_when_ArraySlice_l166_22_2);
  assign _zz_when_ArraySlice_l112_22 = (wReg % _zz__zz_when_ArraySlice_l112_22);
  assign when_ArraySlice_l112_22 = (_zz_when_ArraySlice_l112_22 != 6'h0);
  assign when_ArraySlice_l113_22 = (7'h40 <= _zz_when_ArraySlice_l113_22);
  always @(*) begin
    if(when_ArraySlice_l112_22) begin
      if(when_ArraySlice_l113_22) begin
        _zz_when_ArraySlice_l173_22 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_22 = (_zz__zz_when_ArraySlice_l173_22 - _zz__zz_when_ArraySlice_l173_22_3);
      end
    end else begin
      if(when_ArraySlice_l118_22) begin
        _zz_when_ArraySlice_l173_22 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_22 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_22 = (_zz_when_ArraySlice_l118_22 <= wReg);
  assign when_ArraySlice_l173_22 = (_zz_when_ArraySlice_l173_22_1 <= _zz_when_ArraySlice_l173_22_3);
  assign when_ArraySlice_l165_23 = (_zz_when_ArraySlice_l165_23 <= selectWriteFifo);
  assign when_ArraySlice_l166_23 = (_zz_when_ArraySlice_l166_23 <= _zz_when_ArraySlice_l166_23_2);
  assign _zz_when_ArraySlice_l112_23 = (wReg % _zz__zz_when_ArraySlice_l112_23);
  assign when_ArraySlice_l112_23 = (_zz_when_ArraySlice_l112_23 != 6'h0);
  assign when_ArraySlice_l113_23 = (7'h40 <= _zz_when_ArraySlice_l113_23);
  always @(*) begin
    if(when_ArraySlice_l112_23) begin
      if(when_ArraySlice_l113_23) begin
        _zz_when_ArraySlice_l173_23 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_23 = (_zz__zz_when_ArraySlice_l173_23 - _zz__zz_when_ArraySlice_l173_23_3);
      end
    end else begin
      if(when_ArraySlice_l118_23) begin
        _zz_when_ArraySlice_l173_23 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_23 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_23 = (_zz_when_ArraySlice_l118_23 <= wReg);
  assign when_ArraySlice_l173_23 = (_zz_when_ArraySlice_l173_23_1 <= _zz_when_ArraySlice_l173_23_3);
  assign when_ArraySlice_l418 = (! ((((((_zz_when_ArraySlice_l418 && _zz_when_ArraySlice_l418_1) && (holdReadOp_4 == _zz_when_ArraySlice_l418_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l418_3 && _zz_when_ArraySlice_l418_4) && (debug_4_2 == _zz_when_ArraySlice_l418_5)) && (debug_5_2 == 1'b1)) && (debug_6_2 == 1'b1)) && (debug_7_2 == 1'b1))));
  assign when_ArraySlice_l421 = (wReg <= _zz_when_ArraySlice_l421);
  assign outputStreamArrayData_0_fire_3 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l425 = ((_zz_when_ArraySlice_l425 == 13'h0) && outputStreamArrayData_0_fire_3);
  assign outputStreamArrayData_0_fire_4 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l436 = ((handshakeTimes_0_value == _zz_when_ArraySlice_l436) && outputStreamArrayData_0_fire_4);
  assign _zz_when_ArraySlice_l94_2 = (hReg % _zz__zz_when_ArraySlice_l94_2);
  assign when_ArraySlice_l94_2 = (_zz_when_ArraySlice_l94_2 != 6'h0);
  assign when_ArraySlice_l95_2 = (7'h40 <= _zz_when_ArraySlice_l95_2_1);
  always @(*) begin
    if(when_ArraySlice_l94_2) begin
      if(when_ArraySlice_l95_2) begin
        _zz_when_ArraySlice_l437 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437 = (_zz__zz_when_ArraySlice_l437 - _zz__zz_when_ArraySlice_l437_3);
      end
    end else begin
      if(when_ArraySlice_l99_2) begin
        _zz_when_ArraySlice_l437 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_2 = (_zz_when_ArraySlice_l99_2 <= hReg);
  assign when_ArraySlice_l437 = (_zz_when_ArraySlice_l437_8 < _zz_when_ArraySlice_l437_11);
  always @(*) begin
    debug_0_3 = 1'b0;
    if(when_ArraySlice_l165_24) begin
      if(when_ArraySlice_l166_24) begin
        debug_0_3 = 1'b1;
      end else begin
        debug_0_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_24) begin
        debug_0_3 = 1'b1;
      end else begin
        debug_0_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_3 = 1'b0;
    if(when_ArraySlice_l165_25) begin
      if(when_ArraySlice_l166_25) begin
        debug_1_3 = 1'b1;
      end else begin
        debug_1_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_25) begin
        debug_1_3 = 1'b1;
      end else begin
        debug_1_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_3 = 1'b0;
    if(when_ArraySlice_l165_26) begin
      if(when_ArraySlice_l166_26) begin
        debug_2_3 = 1'b1;
      end else begin
        debug_2_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_26) begin
        debug_2_3 = 1'b1;
      end else begin
        debug_2_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_3 = 1'b0;
    if(when_ArraySlice_l165_27) begin
      if(when_ArraySlice_l166_27) begin
        debug_3_3 = 1'b1;
      end else begin
        debug_3_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_27) begin
        debug_3_3 = 1'b1;
      end else begin
        debug_3_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_3 = 1'b0;
    if(when_ArraySlice_l165_28) begin
      if(when_ArraySlice_l166_28) begin
        debug_4_3 = 1'b1;
      end else begin
        debug_4_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_28) begin
        debug_4_3 = 1'b1;
      end else begin
        debug_4_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_3 = 1'b0;
    if(when_ArraySlice_l165_29) begin
      if(when_ArraySlice_l166_29) begin
        debug_5_3 = 1'b1;
      end else begin
        debug_5_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_29) begin
        debug_5_3 = 1'b1;
      end else begin
        debug_5_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_3 = 1'b0;
    if(when_ArraySlice_l165_30) begin
      if(when_ArraySlice_l166_30) begin
        debug_6_3 = 1'b1;
      end else begin
        debug_6_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_30) begin
        debug_6_3 = 1'b1;
      end else begin
        debug_6_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_3 = 1'b0;
    if(when_ArraySlice_l165_31) begin
      if(when_ArraySlice_l166_31) begin
        debug_7_3 = 1'b1;
      end else begin
        debug_7_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_31) begin
        debug_7_3 = 1'b1;
      end else begin
        debug_7_3 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_24 = (_zz_when_ArraySlice_l165_24 <= selectWriteFifo);
  assign when_ArraySlice_l166_24 = (_zz_when_ArraySlice_l166_24 <= _zz_when_ArraySlice_l166_24_1);
  assign _zz_when_ArraySlice_l112_24 = (wReg % _zz__zz_when_ArraySlice_l112_24);
  assign when_ArraySlice_l112_24 = (_zz_when_ArraySlice_l112_24 != 6'h0);
  assign when_ArraySlice_l113_24 = (7'h40 <= _zz_when_ArraySlice_l113_24);
  always @(*) begin
    if(when_ArraySlice_l112_24) begin
      if(when_ArraySlice_l113_24) begin
        _zz_when_ArraySlice_l173_24 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_24 = (_zz__zz_when_ArraySlice_l173_24 - _zz__zz_when_ArraySlice_l173_24_3);
      end
    end else begin
      if(when_ArraySlice_l118_24) begin
        _zz_when_ArraySlice_l173_24 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_24 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_24 = (_zz_when_ArraySlice_l118_24 <= wReg);
  assign when_ArraySlice_l173_24 = (_zz_when_ArraySlice_l173_24_1 <= _zz_when_ArraySlice_l173_24_2);
  assign when_ArraySlice_l165_25 = (_zz_when_ArraySlice_l165_25 <= selectWriteFifo);
  assign when_ArraySlice_l166_25 = (_zz_when_ArraySlice_l166_25 <= _zz_when_ArraySlice_l166_25_1);
  assign _zz_when_ArraySlice_l112_25 = (wReg % _zz__zz_when_ArraySlice_l112_25);
  assign when_ArraySlice_l112_25 = (_zz_when_ArraySlice_l112_25 != 6'h0);
  assign when_ArraySlice_l113_25 = (7'h40 <= _zz_when_ArraySlice_l113_25);
  always @(*) begin
    if(when_ArraySlice_l112_25) begin
      if(when_ArraySlice_l113_25) begin
        _zz_when_ArraySlice_l173_25 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_25 = (_zz__zz_when_ArraySlice_l173_25 - _zz__zz_when_ArraySlice_l173_25_3);
      end
    end else begin
      if(when_ArraySlice_l118_25) begin
        _zz_when_ArraySlice_l173_25 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_25 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_25 = (_zz_when_ArraySlice_l118_25 <= wReg);
  assign when_ArraySlice_l173_25 = (_zz_when_ArraySlice_l173_25_1 <= _zz_when_ArraySlice_l173_25_3);
  assign when_ArraySlice_l165_26 = (_zz_when_ArraySlice_l165_26 <= selectWriteFifo);
  assign when_ArraySlice_l166_26 = (_zz_when_ArraySlice_l166_26 <= _zz_when_ArraySlice_l166_26_1);
  assign _zz_when_ArraySlice_l112_26 = (wReg % _zz__zz_when_ArraySlice_l112_26);
  assign when_ArraySlice_l112_26 = (_zz_when_ArraySlice_l112_26 != 6'h0);
  assign when_ArraySlice_l113_26 = (7'h40 <= _zz_when_ArraySlice_l113_26);
  always @(*) begin
    if(when_ArraySlice_l112_26) begin
      if(when_ArraySlice_l113_26) begin
        _zz_when_ArraySlice_l173_26 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_26 = (_zz__zz_when_ArraySlice_l173_26 - _zz__zz_when_ArraySlice_l173_26_3);
      end
    end else begin
      if(when_ArraySlice_l118_26) begin
        _zz_when_ArraySlice_l173_26 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_26 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_26 = (_zz_when_ArraySlice_l118_26 <= wReg);
  assign when_ArraySlice_l173_26 = (_zz_when_ArraySlice_l173_26_1 <= _zz_when_ArraySlice_l173_26_3);
  assign when_ArraySlice_l165_27 = (_zz_when_ArraySlice_l165_27 <= selectWriteFifo);
  assign when_ArraySlice_l166_27 = (_zz_when_ArraySlice_l166_27 <= _zz_when_ArraySlice_l166_27_1);
  assign _zz_when_ArraySlice_l112_27 = (wReg % _zz__zz_when_ArraySlice_l112_27);
  assign when_ArraySlice_l112_27 = (_zz_when_ArraySlice_l112_27 != 6'h0);
  assign when_ArraySlice_l113_27 = (7'h40 <= _zz_when_ArraySlice_l113_27);
  always @(*) begin
    if(when_ArraySlice_l112_27) begin
      if(when_ArraySlice_l113_27) begin
        _zz_when_ArraySlice_l173_27 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_27 = (_zz__zz_when_ArraySlice_l173_27 - _zz__zz_when_ArraySlice_l173_27_3);
      end
    end else begin
      if(when_ArraySlice_l118_27) begin
        _zz_when_ArraySlice_l173_27 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_27 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_27 = (_zz_when_ArraySlice_l118_27 <= wReg);
  assign when_ArraySlice_l173_27 = (_zz_when_ArraySlice_l173_27_1 <= _zz_when_ArraySlice_l173_27_3);
  assign when_ArraySlice_l165_28 = (_zz_when_ArraySlice_l165_28 <= selectWriteFifo);
  assign when_ArraySlice_l166_28 = (_zz_when_ArraySlice_l166_28 <= _zz_when_ArraySlice_l166_28_1);
  assign _zz_when_ArraySlice_l112_28 = (wReg % _zz__zz_when_ArraySlice_l112_28);
  assign when_ArraySlice_l112_28 = (_zz_when_ArraySlice_l112_28 != 6'h0);
  assign when_ArraySlice_l113_28 = (7'h40 <= _zz_when_ArraySlice_l113_28);
  always @(*) begin
    if(when_ArraySlice_l112_28) begin
      if(when_ArraySlice_l113_28) begin
        _zz_when_ArraySlice_l173_28 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_28 = (_zz__zz_when_ArraySlice_l173_28 - _zz__zz_when_ArraySlice_l173_28_3);
      end
    end else begin
      if(when_ArraySlice_l118_28) begin
        _zz_when_ArraySlice_l173_28 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_28 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_28 = (_zz_when_ArraySlice_l118_28 <= wReg);
  assign when_ArraySlice_l173_28 = (_zz_when_ArraySlice_l173_28_1 <= _zz_when_ArraySlice_l173_28_3);
  assign when_ArraySlice_l165_29 = (_zz_when_ArraySlice_l165_29 <= selectWriteFifo);
  assign when_ArraySlice_l166_29 = (_zz_when_ArraySlice_l166_29 <= _zz_when_ArraySlice_l166_29_2);
  assign _zz_when_ArraySlice_l112_29 = (wReg % _zz__zz_when_ArraySlice_l112_29);
  assign when_ArraySlice_l112_29 = (_zz_when_ArraySlice_l112_29 != 6'h0);
  assign when_ArraySlice_l113_29 = (7'h40 <= _zz_when_ArraySlice_l113_29);
  always @(*) begin
    if(when_ArraySlice_l112_29) begin
      if(when_ArraySlice_l113_29) begin
        _zz_when_ArraySlice_l173_29 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_29 = (_zz__zz_when_ArraySlice_l173_29 - _zz__zz_when_ArraySlice_l173_29_3);
      end
    end else begin
      if(when_ArraySlice_l118_29) begin
        _zz_when_ArraySlice_l173_29 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_29 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_29 = (_zz_when_ArraySlice_l118_29 <= wReg);
  assign when_ArraySlice_l173_29 = (_zz_when_ArraySlice_l173_29_1 <= _zz_when_ArraySlice_l173_29_3);
  assign when_ArraySlice_l165_30 = (_zz_when_ArraySlice_l165_30 <= selectWriteFifo);
  assign when_ArraySlice_l166_30 = (_zz_when_ArraySlice_l166_30 <= _zz_when_ArraySlice_l166_30_2);
  assign _zz_when_ArraySlice_l112_30 = (wReg % _zz__zz_when_ArraySlice_l112_30);
  assign when_ArraySlice_l112_30 = (_zz_when_ArraySlice_l112_30 != 6'h0);
  assign when_ArraySlice_l113_30 = (7'h40 <= _zz_when_ArraySlice_l113_30);
  always @(*) begin
    if(when_ArraySlice_l112_30) begin
      if(when_ArraySlice_l113_30) begin
        _zz_when_ArraySlice_l173_30 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_30 = (_zz__zz_when_ArraySlice_l173_30 - _zz__zz_when_ArraySlice_l173_30_3);
      end
    end else begin
      if(when_ArraySlice_l118_30) begin
        _zz_when_ArraySlice_l173_30 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_30 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_30 = (_zz_when_ArraySlice_l118_30 <= wReg);
  assign when_ArraySlice_l173_30 = (_zz_when_ArraySlice_l173_30_1 <= _zz_when_ArraySlice_l173_30_3);
  assign when_ArraySlice_l165_31 = (_zz_when_ArraySlice_l165_31 <= selectWriteFifo);
  assign when_ArraySlice_l166_31 = (_zz_when_ArraySlice_l166_31 <= _zz_when_ArraySlice_l166_31_2);
  assign _zz_when_ArraySlice_l112_31 = (wReg % _zz__zz_when_ArraySlice_l112_31);
  assign when_ArraySlice_l112_31 = (_zz_when_ArraySlice_l112_31 != 6'h0);
  assign when_ArraySlice_l113_31 = (7'h40 <= _zz_when_ArraySlice_l113_31);
  always @(*) begin
    if(when_ArraySlice_l112_31) begin
      if(when_ArraySlice_l113_31) begin
        _zz_when_ArraySlice_l173_31 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_31 = (_zz__zz_when_ArraySlice_l173_31 - _zz__zz_when_ArraySlice_l173_31_3);
      end
    end else begin
      if(when_ArraySlice_l118_31) begin
        _zz_when_ArraySlice_l173_31 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_31 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_31 = (_zz_when_ArraySlice_l118_31 <= wReg);
  assign when_ArraySlice_l173_31 = (_zz_when_ArraySlice_l173_31_1 <= _zz_when_ArraySlice_l173_31_3);
  assign when_ArraySlice_l444 = (! ((((((_zz_when_ArraySlice_l444 && _zz_when_ArraySlice_l444_1) && (holdReadOp_4 == _zz_when_ArraySlice_l444_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l444_3 && _zz_when_ArraySlice_l444_4) && (debug_4_3 == _zz_when_ArraySlice_l444_5)) && (debug_5_3 == 1'b1)) && (debug_6_3 == 1'b1)) && (debug_7_3 == 1'b1))));
  assign outputStreamArrayData_0_fire_5 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l448 = ((_zz_when_ArraySlice_l448 == 13'h0) && outputStreamArrayData_0_fire_5);
  assign when_ArraySlice_l434 = (allowPadding_0 && (wReg <= _zz_when_ArraySlice_l434));
  assign outputStreamArrayData_0_fire_6 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l455 = (handshakeTimes_0_value == _zz_when_ArraySlice_l455);
  assign when_ArraySlice_l373_1 = (_zz_when_ArraySlice_l373_1_1 < wReg);
  assign when_ArraySlice_l374_1 = ((! holdReadOp_1) && (_zz_when_ArraySlice_l374_1_1 != 7'h0));
  assign _zz_outputStreamArrayData_1_valid = (selectReadFifo_1 + _zz__zz_outputStreamArrayData_1_valid);
  assign _zz_4 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_1_valid);
  assign _zz_io_pop_ready_1 = outputStreamArrayData_1_ready;
  assign when_ArraySlice_l379_1 = (! holdReadOp_1);
  assign outputStreamArrayData_1_fire = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l380_1 = ((_zz_when_ArraySlice_l380_1_1 < _zz_when_ArraySlice_l380_1_3) && outputStreamArrayData_1_fire);
  assign when_ArraySlice_l381_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l381_1_1);
  assign when_ArraySlice_l384_1 = (_zz_when_ArraySlice_l384_1_1 == 13'h0);
  assign outputStreamArrayData_1_fire_1 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l389_1 = ((_zz_when_ArraySlice_l389_1_1 == _zz_when_ArraySlice_l389_1_5) && outputStreamArrayData_1_fire_1);
  assign when_ArraySlice_l390_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l390_1_1);
  assign _zz_when_ArraySlice_l94_3 = (hReg % _zz__zz_when_ArraySlice_l94_3);
  assign when_ArraySlice_l94_3 = (_zz_when_ArraySlice_l94_3 != 6'h0);
  assign when_ArraySlice_l95_3 = (7'h40 <= _zz_when_ArraySlice_l95_3_1);
  always @(*) begin
    if(when_ArraySlice_l94_3) begin
      if(when_ArraySlice_l95_3) begin
        _zz_when_ArraySlice_l392_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_1 = (_zz__zz_when_ArraySlice_l392_1_1 - _zz__zz_when_ArraySlice_l392_1_4);
      end
    end else begin
      if(when_ArraySlice_l99_3) begin
        _zz_when_ArraySlice_l392_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_1 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_3 = (_zz_when_ArraySlice_l99_3 <= hReg);
  assign when_ArraySlice_l392_1 = (_zz_when_ArraySlice_l392_1_1 < _zz_when_ArraySlice_l392_1_4);
  always @(*) begin
    debug_0_4 = 1'b0;
    if(when_ArraySlice_l165_32) begin
      if(when_ArraySlice_l166_32) begin
        debug_0_4 = 1'b1;
      end else begin
        debug_0_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_32) begin
        debug_0_4 = 1'b1;
      end else begin
        debug_0_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_4 = 1'b0;
    if(when_ArraySlice_l165_33) begin
      if(when_ArraySlice_l166_33) begin
        debug_1_4 = 1'b1;
      end else begin
        debug_1_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_33) begin
        debug_1_4 = 1'b1;
      end else begin
        debug_1_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_4 = 1'b0;
    if(when_ArraySlice_l165_34) begin
      if(when_ArraySlice_l166_34) begin
        debug_2_4 = 1'b1;
      end else begin
        debug_2_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_34) begin
        debug_2_4 = 1'b1;
      end else begin
        debug_2_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_4 = 1'b0;
    if(when_ArraySlice_l165_35) begin
      if(when_ArraySlice_l166_35) begin
        debug_3_4 = 1'b1;
      end else begin
        debug_3_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_35) begin
        debug_3_4 = 1'b1;
      end else begin
        debug_3_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_4 = 1'b0;
    if(when_ArraySlice_l165_36) begin
      if(when_ArraySlice_l166_36) begin
        debug_4_4 = 1'b1;
      end else begin
        debug_4_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_36) begin
        debug_4_4 = 1'b1;
      end else begin
        debug_4_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_4 = 1'b0;
    if(when_ArraySlice_l165_37) begin
      if(when_ArraySlice_l166_37) begin
        debug_5_4 = 1'b1;
      end else begin
        debug_5_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_37) begin
        debug_5_4 = 1'b1;
      end else begin
        debug_5_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_4 = 1'b0;
    if(when_ArraySlice_l165_38) begin
      if(when_ArraySlice_l166_38) begin
        debug_6_4 = 1'b1;
      end else begin
        debug_6_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_38) begin
        debug_6_4 = 1'b1;
      end else begin
        debug_6_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_4 = 1'b0;
    if(when_ArraySlice_l165_39) begin
      if(when_ArraySlice_l166_39) begin
        debug_7_4 = 1'b1;
      end else begin
        debug_7_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_39) begin
        debug_7_4 = 1'b1;
      end else begin
        debug_7_4 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_32 = (_zz_when_ArraySlice_l165_32 <= selectWriteFifo);
  assign when_ArraySlice_l166_32 = (_zz_when_ArraySlice_l166_32 <= _zz_when_ArraySlice_l166_32_1);
  assign _zz_when_ArraySlice_l112_32 = (wReg % _zz__zz_when_ArraySlice_l112_32);
  assign when_ArraySlice_l112_32 = (_zz_when_ArraySlice_l112_32 != 6'h0);
  assign when_ArraySlice_l113_32 = (7'h40 <= _zz_when_ArraySlice_l113_32);
  always @(*) begin
    if(when_ArraySlice_l112_32) begin
      if(when_ArraySlice_l113_32) begin
        _zz_when_ArraySlice_l173_32 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_32 = (_zz__zz_when_ArraySlice_l173_32 - _zz__zz_when_ArraySlice_l173_32_3);
      end
    end else begin
      if(when_ArraySlice_l118_32) begin
        _zz_when_ArraySlice_l173_32 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_32 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_32 = (_zz_when_ArraySlice_l118_32 <= wReg);
  assign when_ArraySlice_l173_32 = (_zz_when_ArraySlice_l173_32_1 <= _zz_when_ArraySlice_l173_32_2);
  assign when_ArraySlice_l165_33 = (_zz_when_ArraySlice_l165_33 <= selectWriteFifo);
  assign when_ArraySlice_l166_33 = (_zz_when_ArraySlice_l166_33 <= _zz_when_ArraySlice_l166_33_1);
  assign _zz_when_ArraySlice_l112_33 = (wReg % _zz__zz_when_ArraySlice_l112_33);
  assign when_ArraySlice_l112_33 = (_zz_when_ArraySlice_l112_33 != 6'h0);
  assign when_ArraySlice_l113_33 = (7'h40 <= _zz_when_ArraySlice_l113_33);
  always @(*) begin
    if(when_ArraySlice_l112_33) begin
      if(when_ArraySlice_l113_33) begin
        _zz_when_ArraySlice_l173_33 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_33 = (_zz__zz_when_ArraySlice_l173_33 - _zz__zz_when_ArraySlice_l173_33_3);
      end
    end else begin
      if(when_ArraySlice_l118_33) begin
        _zz_when_ArraySlice_l173_33 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_33 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_33 = (_zz_when_ArraySlice_l118_33 <= wReg);
  assign when_ArraySlice_l173_33 = (_zz_when_ArraySlice_l173_33_1 <= _zz_when_ArraySlice_l173_33_3);
  assign when_ArraySlice_l165_34 = (_zz_when_ArraySlice_l165_34 <= selectWriteFifo);
  assign when_ArraySlice_l166_34 = (_zz_when_ArraySlice_l166_34 <= _zz_when_ArraySlice_l166_34_1);
  assign _zz_when_ArraySlice_l112_34 = (wReg % _zz__zz_when_ArraySlice_l112_34);
  assign when_ArraySlice_l112_34 = (_zz_when_ArraySlice_l112_34 != 6'h0);
  assign when_ArraySlice_l113_34 = (7'h40 <= _zz_when_ArraySlice_l113_34);
  always @(*) begin
    if(when_ArraySlice_l112_34) begin
      if(when_ArraySlice_l113_34) begin
        _zz_when_ArraySlice_l173_34 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_34 = (_zz__zz_when_ArraySlice_l173_34 - _zz__zz_when_ArraySlice_l173_34_3);
      end
    end else begin
      if(when_ArraySlice_l118_34) begin
        _zz_when_ArraySlice_l173_34 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_34 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_34 = (_zz_when_ArraySlice_l118_34 <= wReg);
  assign when_ArraySlice_l173_34 = (_zz_when_ArraySlice_l173_34_1 <= _zz_when_ArraySlice_l173_34_3);
  assign when_ArraySlice_l165_35 = (_zz_when_ArraySlice_l165_35 <= selectWriteFifo);
  assign when_ArraySlice_l166_35 = (_zz_when_ArraySlice_l166_35 <= _zz_when_ArraySlice_l166_35_1);
  assign _zz_when_ArraySlice_l112_35 = (wReg % _zz__zz_when_ArraySlice_l112_35);
  assign when_ArraySlice_l112_35 = (_zz_when_ArraySlice_l112_35 != 6'h0);
  assign when_ArraySlice_l113_35 = (7'h40 <= _zz_when_ArraySlice_l113_35);
  always @(*) begin
    if(when_ArraySlice_l112_35) begin
      if(when_ArraySlice_l113_35) begin
        _zz_when_ArraySlice_l173_35 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_35 = (_zz__zz_when_ArraySlice_l173_35 - _zz__zz_when_ArraySlice_l173_35_3);
      end
    end else begin
      if(when_ArraySlice_l118_35) begin
        _zz_when_ArraySlice_l173_35 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_35 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_35 = (_zz_when_ArraySlice_l118_35 <= wReg);
  assign when_ArraySlice_l173_35 = (_zz_when_ArraySlice_l173_35_1 <= _zz_when_ArraySlice_l173_35_3);
  assign when_ArraySlice_l165_36 = (_zz_when_ArraySlice_l165_36 <= selectWriteFifo);
  assign when_ArraySlice_l166_36 = (_zz_when_ArraySlice_l166_36 <= _zz_when_ArraySlice_l166_36_1);
  assign _zz_when_ArraySlice_l112_36 = (wReg % _zz__zz_when_ArraySlice_l112_36);
  assign when_ArraySlice_l112_36 = (_zz_when_ArraySlice_l112_36 != 6'h0);
  assign when_ArraySlice_l113_36 = (7'h40 <= _zz_when_ArraySlice_l113_36);
  always @(*) begin
    if(when_ArraySlice_l112_36) begin
      if(when_ArraySlice_l113_36) begin
        _zz_when_ArraySlice_l173_36 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_36 = (_zz__zz_when_ArraySlice_l173_36 - _zz__zz_when_ArraySlice_l173_36_3);
      end
    end else begin
      if(when_ArraySlice_l118_36) begin
        _zz_when_ArraySlice_l173_36 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_36 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_36 = (_zz_when_ArraySlice_l118_36 <= wReg);
  assign when_ArraySlice_l173_36 = (_zz_when_ArraySlice_l173_36_1 <= _zz_when_ArraySlice_l173_36_3);
  assign when_ArraySlice_l165_37 = (_zz_when_ArraySlice_l165_37 <= selectWriteFifo);
  assign when_ArraySlice_l166_37 = (_zz_when_ArraySlice_l166_37 <= _zz_when_ArraySlice_l166_37_2);
  assign _zz_when_ArraySlice_l112_37 = (wReg % _zz__zz_when_ArraySlice_l112_37);
  assign when_ArraySlice_l112_37 = (_zz_when_ArraySlice_l112_37 != 6'h0);
  assign when_ArraySlice_l113_37 = (7'h40 <= _zz_when_ArraySlice_l113_37);
  always @(*) begin
    if(when_ArraySlice_l112_37) begin
      if(when_ArraySlice_l113_37) begin
        _zz_when_ArraySlice_l173_37 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_37 = (_zz__zz_when_ArraySlice_l173_37 - _zz__zz_when_ArraySlice_l173_37_3);
      end
    end else begin
      if(when_ArraySlice_l118_37) begin
        _zz_when_ArraySlice_l173_37 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_37 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_37 = (_zz_when_ArraySlice_l118_37 <= wReg);
  assign when_ArraySlice_l173_37 = (_zz_when_ArraySlice_l173_37_1 <= _zz_when_ArraySlice_l173_37_3);
  assign when_ArraySlice_l165_38 = (_zz_when_ArraySlice_l165_38 <= selectWriteFifo);
  assign when_ArraySlice_l166_38 = (_zz_when_ArraySlice_l166_38 <= _zz_when_ArraySlice_l166_38_2);
  assign _zz_when_ArraySlice_l112_38 = (wReg % _zz__zz_when_ArraySlice_l112_38);
  assign when_ArraySlice_l112_38 = (_zz_when_ArraySlice_l112_38 != 6'h0);
  assign when_ArraySlice_l113_38 = (7'h40 <= _zz_when_ArraySlice_l113_38);
  always @(*) begin
    if(when_ArraySlice_l112_38) begin
      if(when_ArraySlice_l113_38) begin
        _zz_when_ArraySlice_l173_38 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_38 = (_zz__zz_when_ArraySlice_l173_38 - _zz__zz_when_ArraySlice_l173_38_3);
      end
    end else begin
      if(when_ArraySlice_l118_38) begin
        _zz_when_ArraySlice_l173_38 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_38 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_38 = (_zz_when_ArraySlice_l118_38 <= wReg);
  assign when_ArraySlice_l173_38 = (_zz_when_ArraySlice_l173_38_1 <= _zz_when_ArraySlice_l173_38_3);
  assign when_ArraySlice_l165_39 = (_zz_when_ArraySlice_l165_39 <= selectWriteFifo);
  assign when_ArraySlice_l166_39 = (_zz_when_ArraySlice_l166_39 <= _zz_when_ArraySlice_l166_39_2);
  assign _zz_when_ArraySlice_l112_39 = (wReg % _zz__zz_when_ArraySlice_l112_39);
  assign when_ArraySlice_l112_39 = (_zz_when_ArraySlice_l112_39 != 6'h0);
  assign when_ArraySlice_l113_39 = (7'h40 <= _zz_when_ArraySlice_l113_39);
  always @(*) begin
    if(when_ArraySlice_l112_39) begin
      if(when_ArraySlice_l113_39) begin
        _zz_when_ArraySlice_l173_39 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_39 = (_zz__zz_when_ArraySlice_l173_39 - _zz__zz_when_ArraySlice_l173_39_3);
      end
    end else begin
      if(when_ArraySlice_l118_39) begin
        _zz_when_ArraySlice_l173_39 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_39 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_39 = (_zz_when_ArraySlice_l118_39 <= wReg);
  assign when_ArraySlice_l173_39 = (_zz_when_ArraySlice_l173_39_1 <= _zz_when_ArraySlice_l173_39_3);
  assign when_ArraySlice_l398_1 = (! ((((((_zz_when_ArraySlice_l398_1_1 && _zz_when_ArraySlice_l398_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l398_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l398_1_4 && _zz_when_ArraySlice_l398_1_5) && (debug_4_4 == _zz_when_ArraySlice_l398_1_6)) && (debug_5_4 == 1'b1)) && (debug_6_4 == 1'b1)) && (debug_7_4 == 1'b1))));
  assign when_ArraySlice_l401_1 = (wReg <= _zz_when_ArraySlice_l401_1_1);
  assign when_ArraySlice_l405_1 = (_zz_when_ArraySlice_l405_1_1 == 13'h0);
  assign when_ArraySlice_l409_1 = (_zz_when_ArraySlice_l409_1_1 == 7'h0);
  assign outputStreamArrayData_1_fire_2 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l410_1 = ((handshakeTimes_1_value == _zz_when_ArraySlice_l410_1_1) && outputStreamArrayData_1_fire_2);
  assign _zz_when_ArraySlice_l94_4 = (hReg % _zz__zz_when_ArraySlice_l94_4);
  assign when_ArraySlice_l94_4 = (_zz_when_ArraySlice_l94_4 != 6'h0);
  assign when_ArraySlice_l95_4 = (7'h40 <= _zz_when_ArraySlice_l95_4_1);
  always @(*) begin
    if(when_ArraySlice_l94_4) begin
      if(when_ArraySlice_l95_4) begin
        _zz_when_ArraySlice_l412_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_1 = (_zz__zz_when_ArraySlice_l412_1_1 - _zz__zz_when_ArraySlice_l412_1_4);
      end
    end else begin
      if(when_ArraySlice_l99_4) begin
        _zz_when_ArraySlice_l412_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_1 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_4 = (_zz_when_ArraySlice_l99_4 <= hReg);
  assign when_ArraySlice_l412_1 = (_zz_when_ArraySlice_l412_1_1 < _zz_when_ArraySlice_l412_1_4);
  always @(*) begin
    debug_0_5 = 1'b0;
    if(when_ArraySlice_l165_40) begin
      if(when_ArraySlice_l166_40) begin
        debug_0_5 = 1'b1;
      end else begin
        debug_0_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_40) begin
        debug_0_5 = 1'b1;
      end else begin
        debug_0_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_5 = 1'b0;
    if(when_ArraySlice_l165_41) begin
      if(when_ArraySlice_l166_41) begin
        debug_1_5 = 1'b1;
      end else begin
        debug_1_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_41) begin
        debug_1_5 = 1'b1;
      end else begin
        debug_1_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_5 = 1'b0;
    if(when_ArraySlice_l165_42) begin
      if(when_ArraySlice_l166_42) begin
        debug_2_5 = 1'b1;
      end else begin
        debug_2_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_42) begin
        debug_2_5 = 1'b1;
      end else begin
        debug_2_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_5 = 1'b0;
    if(when_ArraySlice_l165_43) begin
      if(when_ArraySlice_l166_43) begin
        debug_3_5 = 1'b1;
      end else begin
        debug_3_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_43) begin
        debug_3_5 = 1'b1;
      end else begin
        debug_3_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_5 = 1'b0;
    if(when_ArraySlice_l165_44) begin
      if(when_ArraySlice_l166_44) begin
        debug_4_5 = 1'b1;
      end else begin
        debug_4_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_44) begin
        debug_4_5 = 1'b1;
      end else begin
        debug_4_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_5 = 1'b0;
    if(when_ArraySlice_l165_45) begin
      if(when_ArraySlice_l166_45) begin
        debug_5_5 = 1'b1;
      end else begin
        debug_5_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_45) begin
        debug_5_5 = 1'b1;
      end else begin
        debug_5_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_5 = 1'b0;
    if(when_ArraySlice_l165_46) begin
      if(when_ArraySlice_l166_46) begin
        debug_6_5 = 1'b1;
      end else begin
        debug_6_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_46) begin
        debug_6_5 = 1'b1;
      end else begin
        debug_6_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_5 = 1'b0;
    if(when_ArraySlice_l165_47) begin
      if(when_ArraySlice_l166_47) begin
        debug_7_5 = 1'b1;
      end else begin
        debug_7_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_47) begin
        debug_7_5 = 1'b1;
      end else begin
        debug_7_5 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_40 = (_zz_when_ArraySlice_l165_40 <= selectWriteFifo);
  assign when_ArraySlice_l166_40 = (_zz_when_ArraySlice_l166_40 <= _zz_when_ArraySlice_l166_40_1);
  assign _zz_when_ArraySlice_l112_40 = (wReg % _zz__zz_when_ArraySlice_l112_40);
  assign when_ArraySlice_l112_40 = (_zz_when_ArraySlice_l112_40 != 6'h0);
  assign when_ArraySlice_l113_40 = (7'h40 <= _zz_when_ArraySlice_l113_40);
  always @(*) begin
    if(when_ArraySlice_l112_40) begin
      if(when_ArraySlice_l113_40) begin
        _zz_when_ArraySlice_l173_40 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_40 = (_zz__zz_when_ArraySlice_l173_40 - _zz__zz_when_ArraySlice_l173_40_3);
      end
    end else begin
      if(when_ArraySlice_l118_40) begin
        _zz_when_ArraySlice_l173_40 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_40 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_40 = (_zz_when_ArraySlice_l118_40 <= wReg);
  assign when_ArraySlice_l173_40 = (_zz_when_ArraySlice_l173_40_1 <= _zz_when_ArraySlice_l173_40_2);
  assign when_ArraySlice_l165_41 = (_zz_when_ArraySlice_l165_41 <= selectWriteFifo);
  assign when_ArraySlice_l166_41 = (_zz_when_ArraySlice_l166_41 <= _zz_when_ArraySlice_l166_41_1);
  assign _zz_when_ArraySlice_l112_41 = (wReg % _zz__zz_when_ArraySlice_l112_41);
  assign when_ArraySlice_l112_41 = (_zz_when_ArraySlice_l112_41 != 6'h0);
  assign when_ArraySlice_l113_41 = (7'h40 <= _zz_when_ArraySlice_l113_41);
  always @(*) begin
    if(when_ArraySlice_l112_41) begin
      if(when_ArraySlice_l113_41) begin
        _zz_when_ArraySlice_l173_41 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_41 = (_zz__zz_when_ArraySlice_l173_41 - _zz__zz_when_ArraySlice_l173_41_3);
      end
    end else begin
      if(when_ArraySlice_l118_41) begin
        _zz_when_ArraySlice_l173_41 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_41 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_41 = (_zz_when_ArraySlice_l118_41 <= wReg);
  assign when_ArraySlice_l173_41 = (_zz_when_ArraySlice_l173_41_1 <= _zz_when_ArraySlice_l173_41_3);
  assign when_ArraySlice_l165_42 = (_zz_when_ArraySlice_l165_42 <= selectWriteFifo);
  assign when_ArraySlice_l166_42 = (_zz_when_ArraySlice_l166_42 <= _zz_when_ArraySlice_l166_42_1);
  assign _zz_when_ArraySlice_l112_42 = (wReg % _zz__zz_when_ArraySlice_l112_42);
  assign when_ArraySlice_l112_42 = (_zz_when_ArraySlice_l112_42 != 6'h0);
  assign when_ArraySlice_l113_42 = (7'h40 <= _zz_when_ArraySlice_l113_42);
  always @(*) begin
    if(when_ArraySlice_l112_42) begin
      if(when_ArraySlice_l113_42) begin
        _zz_when_ArraySlice_l173_42 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_42 = (_zz__zz_when_ArraySlice_l173_42 - _zz__zz_when_ArraySlice_l173_42_3);
      end
    end else begin
      if(when_ArraySlice_l118_42) begin
        _zz_when_ArraySlice_l173_42 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_42 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_42 = (_zz_when_ArraySlice_l118_42 <= wReg);
  assign when_ArraySlice_l173_42 = (_zz_when_ArraySlice_l173_42_1 <= _zz_when_ArraySlice_l173_42_3);
  assign when_ArraySlice_l165_43 = (_zz_when_ArraySlice_l165_43 <= selectWriteFifo);
  assign when_ArraySlice_l166_43 = (_zz_when_ArraySlice_l166_43 <= _zz_when_ArraySlice_l166_43_1);
  assign _zz_when_ArraySlice_l112_43 = (wReg % _zz__zz_when_ArraySlice_l112_43);
  assign when_ArraySlice_l112_43 = (_zz_when_ArraySlice_l112_43 != 6'h0);
  assign when_ArraySlice_l113_43 = (7'h40 <= _zz_when_ArraySlice_l113_43);
  always @(*) begin
    if(when_ArraySlice_l112_43) begin
      if(when_ArraySlice_l113_43) begin
        _zz_when_ArraySlice_l173_43 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_43 = (_zz__zz_when_ArraySlice_l173_43 - _zz__zz_when_ArraySlice_l173_43_3);
      end
    end else begin
      if(when_ArraySlice_l118_43) begin
        _zz_when_ArraySlice_l173_43 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_43 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_43 = (_zz_when_ArraySlice_l118_43 <= wReg);
  assign when_ArraySlice_l173_43 = (_zz_when_ArraySlice_l173_43_1 <= _zz_when_ArraySlice_l173_43_3);
  assign when_ArraySlice_l165_44 = (_zz_when_ArraySlice_l165_44 <= selectWriteFifo);
  assign when_ArraySlice_l166_44 = (_zz_when_ArraySlice_l166_44 <= _zz_when_ArraySlice_l166_44_1);
  assign _zz_when_ArraySlice_l112_44 = (wReg % _zz__zz_when_ArraySlice_l112_44);
  assign when_ArraySlice_l112_44 = (_zz_when_ArraySlice_l112_44 != 6'h0);
  assign when_ArraySlice_l113_44 = (7'h40 <= _zz_when_ArraySlice_l113_44);
  always @(*) begin
    if(when_ArraySlice_l112_44) begin
      if(when_ArraySlice_l113_44) begin
        _zz_when_ArraySlice_l173_44 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_44 = (_zz__zz_when_ArraySlice_l173_44 - _zz__zz_when_ArraySlice_l173_44_3);
      end
    end else begin
      if(when_ArraySlice_l118_44) begin
        _zz_when_ArraySlice_l173_44 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_44 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_44 = (_zz_when_ArraySlice_l118_44 <= wReg);
  assign when_ArraySlice_l173_44 = (_zz_when_ArraySlice_l173_44_1 <= _zz_when_ArraySlice_l173_44_3);
  assign when_ArraySlice_l165_45 = (_zz_when_ArraySlice_l165_45 <= selectWriteFifo);
  assign when_ArraySlice_l166_45 = (_zz_when_ArraySlice_l166_45 <= _zz_when_ArraySlice_l166_45_2);
  assign _zz_when_ArraySlice_l112_45 = (wReg % _zz__zz_when_ArraySlice_l112_45);
  assign when_ArraySlice_l112_45 = (_zz_when_ArraySlice_l112_45 != 6'h0);
  assign when_ArraySlice_l113_45 = (7'h40 <= _zz_when_ArraySlice_l113_45);
  always @(*) begin
    if(when_ArraySlice_l112_45) begin
      if(when_ArraySlice_l113_45) begin
        _zz_when_ArraySlice_l173_45 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_45 = (_zz__zz_when_ArraySlice_l173_45 - _zz__zz_when_ArraySlice_l173_45_3);
      end
    end else begin
      if(when_ArraySlice_l118_45) begin
        _zz_when_ArraySlice_l173_45 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_45 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_45 = (_zz_when_ArraySlice_l118_45 <= wReg);
  assign when_ArraySlice_l173_45 = (_zz_when_ArraySlice_l173_45_1 <= _zz_when_ArraySlice_l173_45_3);
  assign when_ArraySlice_l165_46 = (_zz_when_ArraySlice_l165_46 <= selectWriteFifo);
  assign when_ArraySlice_l166_46 = (_zz_when_ArraySlice_l166_46 <= _zz_when_ArraySlice_l166_46_2);
  assign _zz_when_ArraySlice_l112_46 = (wReg % _zz__zz_when_ArraySlice_l112_46);
  assign when_ArraySlice_l112_46 = (_zz_when_ArraySlice_l112_46 != 6'h0);
  assign when_ArraySlice_l113_46 = (7'h40 <= _zz_when_ArraySlice_l113_46);
  always @(*) begin
    if(when_ArraySlice_l112_46) begin
      if(when_ArraySlice_l113_46) begin
        _zz_when_ArraySlice_l173_46 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_46 = (_zz__zz_when_ArraySlice_l173_46 - _zz__zz_when_ArraySlice_l173_46_3);
      end
    end else begin
      if(when_ArraySlice_l118_46) begin
        _zz_when_ArraySlice_l173_46 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_46 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_46 = (_zz_when_ArraySlice_l118_46 <= wReg);
  assign when_ArraySlice_l173_46 = (_zz_when_ArraySlice_l173_46_1 <= _zz_when_ArraySlice_l173_46_3);
  assign when_ArraySlice_l165_47 = (_zz_when_ArraySlice_l165_47 <= selectWriteFifo);
  assign when_ArraySlice_l166_47 = (_zz_when_ArraySlice_l166_47 <= _zz_when_ArraySlice_l166_47_2);
  assign _zz_when_ArraySlice_l112_47 = (wReg % _zz__zz_when_ArraySlice_l112_47);
  assign when_ArraySlice_l112_47 = (_zz_when_ArraySlice_l112_47 != 6'h0);
  assign when_ArraySlice_l113_47 = (7'h40 <= _zz_when_ArraySlice_l113_47);
  always @(*) begin
    if(when_ArraySlice_l112_47) begin
      if(when_ArraySlice_l113_47) begin
        _zz_when_ArraySlice_l173_47 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_47 = (_zz__zz_when_ArraySlice_l173_47 - _zz__zz_when_ArraySlice_l173_47_3);
      end
    end else begin
      if(when_ArraySlice_l118_47) begin
        _zz_when_ArraySlice_l173_47 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_47 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_47 = (_zz_when_ArraySlice_l118_47 <= wReg);
  assign when_ArraySlice_l173_47 = (_zz_when_ArraySlice_l173_47_1 <= _zz_when_ArraySlice_l173_47_3);
  assign when_ArraySlice_l418_1 = (! ((((((_zz_when_ArraySlice_l418_1_1 && _zz_when_ArraySlice_l418_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l418_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l418_1_4 && _zz_when_ArraySlice_l418_1_5) && (debug_4_5 == _zz_when_ArraySlice_l418_1_6)) && (debug_5_5 == 1'b1)) && (debug_6_5 == 1'b1)) && (debug_7_5 == 1'b1))));
  assign when_ArraySlice_l421_1 = (wReg <= _zz_when_ArraySlice_l421_1_1);
  assign outputStreamArrayData_1_fire_3 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l425_1 = ((_zz_when_ArraySlice_l425_1_1 == 13'h0) && outputStreamArrayData_1_fire_3);
  assign outputStreamArrayData_1_fire_4 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l436_1 = ((handshakeTimes_1_value == _zz_when_ArraySlice_l436_1_1) && outputStreamArrayData_1_fire_4);
  assign _zz_when_ArraySlice_l94_5 = (hReg % _zz__zz_when_ArraySlice_l94_5);
  assign when_ArraySlice_l94_5 = (_zz_when_ArraySlice_l94_5 != 6'h0);
  assign when_ArraySlice_l95_5 = (7'h40 <= _zz_when_ArraySlice_l95_5);
  always @(*) begin
    if(when_ArraySlice_l94_5) begin
      if(when_ArraySlice_l95_5) begin
        _zz_when_ArraySlice_l437_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_1 = (_zz__zz_when_ArraySlice_l437_1_1 - _zz__zz_when_ArraySlice_l437_1_4);
      end
    end else begin
      if(when_ArraySlice_l99_5) begin
        _zz_when_ArraySlice_l437_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_1 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_5 = (_zz_when_ArraySlice_l99_5 <= hReg);
  assign when_ArraySlice_l437_1 = (_zz_when_ArraySlice_l437_1_1 < _zz_when_ArraySlice_l437_1_4);
  always @(*) begin
    debug_0_6 = 1'b0;
    if(when_ArraySlice_l165_48) begin
      if(when_ArraySlice_l166_48) begin
        debug_0_6 = 1'b1;
      end else begin
        debug_0_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_48) begin
        debug_0_6 = 1'b1;
      end else begin
        debug_0_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_6 = 1'b0;
    if(when_ArraySlice_l165_49) begin
      if(when_ArraySlice_l166_49) begin
        debug_1_6 = 1'b1;
      end else begin
        debug_1_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_49) begin
        debug_1_6 = 1'b1;
      end else begin
        debug_1_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_6 = 1'b0;
    if(when_ArraySlice_l165_50) begin
      if(when_ArraySlice_l166_50) begin
        debug_2_6 = 1'b1;
      end else begin
        debug_2_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_50) begin
        debug_2_6 = 1'b1;
      end else begin
        debug_2_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_6 = 1'b0;
    if(when_ArraySlice_l165_51) begin
      if(when_ArraySlice_l166_51) begin
        debug_3_6 = 1'b1;
      end else begin
        debug_3_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_51) begin
        debug_3_6 = 1'b1;
      end else begin
        debug_3_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_6 = 1'b0;
    if(when_ArraySlice_l165_52) begin
      if(when_ArraySlice_l166_52) begin
        debug_4_6 = 1'b1;
      end else begin
        debug_4_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_52) begin
        debug_4_6 = 1'b1;
      end else begin
        debug_4_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_6 = 1'b0;
    if(when_ArraySlice_l165_53) begin
      if(when_ArraySlice_l166_53) begin
        debug_5_6 = 1'b1;
      end else begin
        debug_5_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_53) begin
        debug_5_6 = 1'b1;
      end else begin
        debug_5_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_6 = 1'b0;
    if(when_ArraySlice_l165_54) begin
      if(when_ArraySlice_l166_54) begin
        debug_6_6 = 1'b1;
      end else begin
        debug_6_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_54) begin
        debug_6_6 = 1'b1;
      end else begin
        debug_6_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_6 = 1'b0;
    if(when_ArraySlice_l165_55) begin
      if(when_ArraySlice_l166_55) begin
        debug_7_6 = 1'b1;
      end else begin
        debug_7_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_55) begin
        debug_7_6 = 1'b1;
      end else begin
        debug_7_6 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_48 = (_zz_when_ArraySlice_l165_48 <= selectWriteFifo);
  assign when_ArraySlice_l166_48 = (_zz_when_ArraySlice_l166_48 <= _zz_when_ArraySlice_l166_48_1);
  assign _zz_when_ArraySlice_l112_48 = (wReg % _zz__zz_when_ArraySlice_l112_48);
  assign when_ArraySlice_l112_48 = (_zz_when_ArraySlice_l112_48 != 6'h0);
  assign when_ArraySlice_l113_48 = (7'h40 <= _zz_when_ArraySlice_l113_48);
  always @(*) begin
    if(when_ArraySlice_l112_48) begin
      if(when_ArraySlice_l113_48) begin
        _zz_when_ArraySlice_l173_48 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_48 = (_zz__zz_when_ArraySlice_l173_48 - _zz__zz_when_ArraySlice_l173_48_3);
      end
    end else begin
      if(when_ArraySlice_l118_48) begin
        _zz_when_ArraySlice_l173_48 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_48 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_48 = (_zz_when_ArraySlice_l118_48 <= wReg);
  assign when_ArraySlice_l173_48 = (_zz_when_ArraySlice_l173_48_1 <= _zz_when_ArraySlice_l173_48_2);
  assign when_ArraySlice_l165_49 = (_zz_when_ArraySlice_l165_49 <= selectWriteFifo);
  assign when_ArraySlice_l166_49 = (_zz_when_ArraySlice_l166_49 <= _zz_when_ArraySlice_l166_49_1);
  assign _zz_when_ArraySlice_l112_49 = (wReg % _zz__zz_when_ArraySlice_l112_49);
  assign when_ArraySlice_l112_49 = (_zz_when_ArraySlice_l112_49 != 6'h0);
  assign when_ArraySlice_l113_49 = (7'h40 <= _zz_when_ArraySlice_l113_49);
  always @(*) begin
    if(when_ArraySlice_l112_49) begin
      if(when_ArraySlice_l113_49) begin
        _zz_when_ArraySlice_l173_49 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_49 = (_zz__zz_when_ArraySlice_l173_49 - _zz__zz_when_ArraySlice_l173_49_3);
      end
    end else begin
      if(when_ArraySlice_l118_49) begin
        _zz_when_ArraySlice_l173_49 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_49 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_49 = (_zz_when_ArraySlice_l118_49 <= wReg);
  assign when_ArraySlice_l173_49 = (_zz_when_ArraySlice_l173_49_1 <= _zz_when_ArraySlice_l173_49_3);
  assign when_ArraySlice_l165_50 = (_zz_when_ArraySlice_l165_50 <= selectWriteFifo);
  assign when_ArraySlice_l166_50 = (_zz_when_ArraySlice_l166_50 <= _zz_when_ArraySlice_l166_50_1);
  assign _zz_when_ArraySlice_l112_50 = (wReg % _zz__zz_when_ArraySlice_l112_50);
  assign when_ArraySlice_l112_50 = (_zz_when_ArraySlice_l112_50 != 6'h0);
  assign when_ArraySlice_l113_50 = (7'h40 <= _zz_when_ArraySlice_l113_50);
  always @(*) begin
    if(when_ArraySlice_l112_50) begin
      if(when_ArraySlice_l113_50) begin
        _zz_when_ArraySlice_l173_50 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_50 = (_zz__zz_when_ArraySlice_l173_50 - _zz__zz_when_ArraySlice_l173_50_3);
      end
    end else begin
      if(when_ArraySlice_l118_50) begin
        _zz_when_ArraySlice_l173_50 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_50 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_50 = (_zz_when_ArraySlice_l118_50 <= wReg);
  assign when_ArraySlice_l173_50 = (_zz_when_ArraySlice_l173_50_1 <= _zz_when_ArraySlice_l173_50_3);
  assign when_ArraySlice_l165_51 = (_zz_when_ArraySlice_l165_51 <= selectWriteFifo);
  assign when_ArraySlice_l166_51 = (_zz_when_ArraySlice_l166_51 <= _zz_when_ArraySlice_l166_51_1);
  assign _zz_when_ArraySlice_l112_51 = (wReg % _zz__zz_when_ArraySlice_l112_51);
  assign when_ArraySlice_l112_51 = (_zz_when_ArraySlice_l112_51 != 6'h0);
  assign when_ArraySlice_l113_51 = (7'h40 <= _zz_when_ArraySlice_l113_51);
  always @(*) begin
    if(when_ArraySlice_l112_51) begin
      if(when_ArraySlice_l113_51) begin
        _zz_when_ArraySlice_l173_51 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_51 = (_zz__zz_when_ArraySlice_l173_51 - _zz__zz_when_ArraySlice_l173_51_3);
      end
    end else begin
      if(when_ArraySlice_l118_51) begin
        _zz_when_ArraySlice_l173_51 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_51 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_51 = (_zz_when_ArraySlice_l118_51 <= wReg);
  assign when_ArraySlice_l173_51 = (_zz_when_ArraySlice_l173_51_1 <= _zz_when_ArraySlice_l173_51_3);
  assign when_ArraySlice_l165_52 = (_zz_when_ArraySlice_l165_52 <= selectWriteFifo);
  assign when_ArraySlice_l166_52 = (_zz_when_ArraySlice_l166_52 <= _zz_when_ArraySlice_l166_52_1);
  assign _zz_when_ArraySlice_l112_52 = (wReg % _zz__zz_when_ArraySlice_l112_52);
  assign when_ArraySlice_l112_52 = (_zz_when_ArraySlice_l112_52 != 6'h0);
  assign when_ArraySlice_l113_52 = (7'h40 <= _zz_when_ArraySlice_l113_52);
  always @(*) begin
    if(when_ArraySlice_l112_52) begin
      if(when_ArraySlice_l113_52) begin
        _zz_when_ArraySlice_l173_52 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_52 = (_zz__zz_when_ArraySlice_l173_52 - _zz__zz_when_ArraySlice_l173_52_3);
      end
    end else begin
      if(when_ArraySlice_l118_52) begin
        _zz_when_ArraySlice_l173_52 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_52 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_52 = (_zz_when_ArraySlice_l118_52 <= wReg);
  assign when_ArraySlice_l173_52 = (_zz_when_ArraySlice_l173_52_1 <= _zz_when_ArraySlice_l173_52_3);
  assign when_ArraySlice_l165_53 = (_zz_when_ArraySlice_l165_53 <= selectWriteFifo);
  assign when_ArraySlice_l166_53 = (_zz_when_ArraySlice_l166_53 <= _zz_when_ArraySlice_l166_53_2);
  assign _zz_when_ArraySlice_l112_53 = (wReg % _zz__zz_when_ArraySlice_l112_53);
  assign when_ArraySlice_l112_53 = (_zz_when_ArraySlice_l112_53 != 6'h0);
  assign when_ArraySlice_l113_53 = (7'h40 <= _zz_when_ArraySlice_l113_53);
  always @(*) begin
    if(when_ArraySlice_l112_53) begin
      if(when_ArraySlice_l113_53) begin
        _zz_when_ArraySlice_l173_53 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_53 = (_zz__zz_when_ArraySlice_l173_53 - _zz__zz_when_ArraySlice_l173_53_3);
      end
    end else begin
      if(when_ArraySlice_l118_53) begin
        _zz_when_ArraySlice_l173_53 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_53 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_53 = (_zz_when_ArraySlice_l118_53 <= wReg);
  assign when_ArraySlice_l173_53 = (_zz_when_ArraySlice_l173_53_1 <= _zz_when_ArraySlice_l173_53_3);
  assign when_ArraySlice_l165_54 = (_zz_when_ArraySlice_l165_54 <= selectWriteFifo);
  assign when_ArraySlice_l166_54 = (_zz_when_ArraySlice_l166_54 <= _zz_when_ArraySlice_l166_54_2);
  assign _zz_when_ArraySlice_l112_54 = (wReg % _zz__zz_when_ArraySlice_l112_54);
  assign when_ArraySlice_l112_54 = (_zz_when_ArraySlice_l112_54 != 6'h0);
  assign when_ArraySlice_l113_54 = (7'h40 <= _zz_when_ArraySlice_l113_54);
  always @(*) begin
    if(when_ArraySlice_l112_54) begin
      if(when_ArraySlice_l113_54) begin
        _zz_when_ArraySlice_l173_54 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_54 = (_zz__zz_when_ArraySlice_l173_54 - _zz__zz_when_ArraySlice_l173_54_3);
      end
    end else begin
      if(when_ArraySlice_l118_54) begin
        _zz_when_ArraySlice_l173_54 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_54 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_54 = (_zz_when_ArraySlice_l118_54 <= wReg);
  assign when_ArraySlice_l173_54 = (_zz_when_ArraySlice_l173_54_1 <= _zz_when_ArraySlice_l173_54_3);
  assign when_ArraySlice_l165_55 = (_zz_when_ArraySlice_l165_55 <= selectWriteFifo);
  assign when_ArraySlice_l166_55 = (_zz_when_ArraySlice_l166_55 <= _zz_when_ArraySlice_l166_55_2);
  assign _zz_when_ArraySlice_l112_55 = (wReg % _zz__zz_when_ArraySlice_l112_55);
  assign when_ArraySlice_l112_55 = (_zz_when_ArraySlice_l112_55 != 6'h0);
  assign when_ArraySlice_l113_55 = (7'h40 <= _zz_when_ArraySlice_l113_55);
  always @(*) begin
    if(when_ArraySlice_l112_55) begin
      if(when_ArraySlice_l113_55) begin
        _zz_when_ArraySlice_l173_55 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_55 = (_zz__zz_when_ArraySlice_l173_55 - _zz__zz_when_ArraySlice_l173_55_3);
      end
    end else begin
      if(when_ArraySlice_l118_55) begin
        _zz_when_ArraySlice_l173_55 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_55 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_55 = (_zz_when_ArraySlice_l118_55 <= wReg);
  assign when_ArraySlice_l173_55 = (_zz_when_ArraySlice_l173_55_1 <= _zz_when_ArraySlice_l173_55_3);
  assign when_ArraySlice_l444_1 = (! ((((((_zz_when_ArraySlice_l444_1_1 && _zz_when_ArraySlice_l444_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l444_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l444_1_4 && _zz_when_ArraySlice_l444_1_5) && (debug_4_6 == _zz_when_ArraySlice_l444_1_6)) && (debug_5_6 == 1'b1)) && (debug_6_6 == 1'b1)) && (debug_7_6 == 1'b1))));
  assign outputStreamArrayData_1_fire_5 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l448_1 = ((_zz_when_ArraySlice_l448_1_1 == 13'h0) && outputStreamArrayData_1_fire_5);
  assign when_ArraySlice_l434_1 = (allowPadding_1 && (wReg <= _zz_when_ArraySlice_l434_1_1));
  assign outputStreamArrayData_1_fire_6 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l455_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l455_1_1);
  assign when_ArraySlice_l373_2 = (_zz_when_ArraySlice_l373_2_1 < wReg);
  assign when_ArraySlice_l374_2 = ((! holdReadOp_2) && (_zz_when_ArraySlice_l374_2_1 != 7'h0));
  assign _zz_outputStreamArrayData_2_valid = (selectReadFifo_2 + _zz__zz_outputStreamArrayData_2_valid);
  assign _zz_5 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_2_valid);
  assign _zz_io_pop_ready_2 = outputStreamArrayData_2_ready;
  assign when_ArraySlice_l379_2 = (! holdReadOp_2);
  assign outputStreamArrayData_2_fire = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l380_2 = ((_zz_when_ArraySlice_l380_2_1 < _zz_when_ArraySlice_l380_2_3) && outputStreamArrayData_2_fire);
  assign when_ArraySlice_l381_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l381_2_1);
  assign when_ArraySlice_l384_2 = (_zz_when_ArraySlice_l384_2_1 == 13'h0);
  assign outputStreamArrayData_2_fire_1 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l389_2 = ((_zz_when_ArraySlice_l389_2_1 == _zz_when_ArraySlice_l389_2_5) && outputStreamArrayData_2_fire_1);
  assign when_ArraySlice_l390_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l390_2_1);
  assign _zz_when_ArraySlice_l94_6 = (hReg % _zz__zz_when_ArraySlice_l94_6);
  assign when_ArraySlice_l94_6 = (_zz_when_ArraySlice_l94_6 != 6'h0);
  assign when_ArraySlice_l95_6 = (7'h40 <= _zz_when_ArraySlice_l95_6);
  always @(*) begin
    if(when_ArraySlice_l94_6) begin
      if(when_ArraySlice_l95_6) begin
        _zz_when_ArraySlice_l392_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_2 = (_zz__zz_when_ArraySlice_l392_2_1 - _zz__zz_when_ArraySlice_l392_2_4);
      end
    end else begin
      if(when_ArraySlice_l99_6) begin
        _zz_when_ArraySlice_l392_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_2 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_6 = (_zz_when_ArraySlice_l99_6 <= hReg);
  assign when_ArraySlice_l392_2 = (_zz_when_ArraySlice_l392_2_1 < _zz_when_ArraySlice_l392_2_4);
  always @(*) begin
    debug_0_7 = 1'b0;
    if(when_ArraySlice_l165_56) begin
      if(when_ArraySlice_l166_56) begin
        debug_0_7 = 1'b1;
      end else begin
        debug_0_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_56) begin
        debug_0_7 = 1'b1;
      end else begin
        debug_0_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_7 = 1'b0;
    if(when_ArraySlice_l165_57) begin
      if(when_ArraySlice_l166_57) begin
        debug_1_7 = 1'b1;
      end else begin
        debug_1_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_57) begin
        debug_1_7 = 1'b1;
      end else begin
        debug_1_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_7 = 1'b0;
    if(when_ArraySlice_l165_58) begin
      if(when_ArraySlice_l166_58) begin
        debug_2_7 = 1'b1;
      end else begin
        debug_2_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_58) begin
        debug_2_7 = 1'b1;
      end else begin
        debug_2_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_7 = 1'b0;
    if(when_ArraySlice_l165_59) begin
      if(when_ArraySlice_l166_59) begin
        debug_3_7 = 1'b1;
      end else begin
        debug_3_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_59) begin
        debug_3_7 = 1'b1;
      end else begin
        debug_3_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_7 = 1'b0;
    if(when_ArraySlice_l165_60) begin
      if(when_ArraySlice_l166_60) begin
        debug_4_7 = 1'b1;
      end else begin
        debug_4_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_60) begin
        debug_4_7 = 1'b1;
      end else begin
        debug_4_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_7 = 1'b0;
    if(when_ArraySlice_l165_61) begin
      if(when_ArraySlice_l166_61) begin
        debug_5_7 = 1'b1;
      end else begin
        debug_5_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_61) begin
        debug_5_7 = 1'b1;
      end else begin
        debug_5_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_7 = 1'b0;
    if(when_ArraySlice_l165_62) begin
      if(when_ArraySlice_l166_62) begin
        debug_6_7 = 1'b1;
      end else begin
        debug_6_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_62) begin
        debug_6_7 = 1'b1;
      end else begin
        debug_6_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_7 = 1'b0;
    if(when_ArraySlice_l165_63) begin
      if(when_ArraySlice_l166_63) begin
        debug_7_7 = 1'b1;
      end else begin
        debug_7_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_63) begin
        debug_7_7 = 1'b1;
      end else begin
        debug_7_7 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_56 = (_zz_when_ArraySlice_l165_56 <= selectWriteFifo);
  assign when_ArraySlice_l166_56 = (_zz_when_ArraySlice_l166_56 <= _zz_when_ArraySlice_l166_56_1);
  assign _zz_when_ArraySlice_l112_56 = (wReg % _zz__zz_when_ArraySlice_l112_56);
  assign when_ArraySlice_l112_56 = (_zz_when_ArraySlice_l112_56 != 6'h0);
  assign when_ArraySlice_l113_56 = (7'h40 <= _zz_when_ArraySlice_l113_56);
  always @(*) begin
    if(when_ArraySlice_l112_56) begin
      if(when_ArraySlice_l113_56) begin
        _zz_when_ArraySlice_l173_56 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_56 = (_zz__zz_when_ArraySlice_l173_56 - _zz__zz_when_ArraySlice_l173_56_3);
      end
    end else begin
      if(when_ArraySlice_l118_56) begin
        _zz_when_ArraySlice_l173_56 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_56 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_56 = (_zz_when_ArraySlice_l118_56 <= wReg);
  assign when_ArraySlice_l173_56 = (_zz_when_ArraySlice_l173_56_1 <= _zz_when_ArraySlice_l173_56_2);
  assign when_ArraySlice_l165_57 = (_zz_when_ArraySlice_l165_57 <= selectWriteFifo);
  assign when_ArraySlice_l166_57 = (_zz_when_ArraySlice_l166_57 <= _zz_when_ArraySlice_l166_57_1);
  assign _zz_when_ArraySlice_l112_57 = (wReg % _zz__zz_when_ArraySlice_l112_57);
  assign when_ArraySlice_l112_57 = (_zz_when_ArraySlice_l112_57 != 6'h0);
  assign when_ArraySlice_l113_57 = (7'h40 <= _zz_when_ArraySlice_l113_57);
  always @(*) begin
    if(when_ArraySlice_l112_57) begin
      if(when_ArraySlice_l113_57) begin
        _zz_when_ArraySlice_l173_57 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_57 = (_zz__zz_when_ArraySlice_l173_57 - _zz__zz_when_ArraySlice_l173_57_3);
      end
    end else begin
      if(when_ArraySlice_l118_57) begin
        _zz_when_ArraySlice_l173_57 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_57 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_57 = (_zz_when_ArraySlice_l118_57 <= wReg);
  assign when_ArraySlice_l173_57 = (_zz_when_ArraySlice_l173_57_1 <= _zz_when_ArraySlice_l173_57_3);
  assign when_ArraySlice_l165_58 = (_zz_when_ArraySlice_l165_58 <= selectWriteFifo);
  assign when_ArraySlice_l166_58 = (_zz_when_ArraySlice_l166_58 <= _zz_when_ArraySlice_l166_58_1);
  assign _zz_when_ArraySlice_l112_58 = (wReg % _zz__zz_when_ArraySlice_l112_58);
  assign when_ArraySlice_l112_58 = (_zz_when_ArraySlice_l112_58 != 6'h0);
  assign when_ArraySlice_l113_58 = (7'h40 <= _zz_when_ArraySlice_l113_58);
  always @(*) begin
    if(when_ArraySlice_l112_58) begin
      if(when_ArraySlice_l113_58) begin
        _zz_when_ArraySlice_l173_58 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_58 = (_zz__zz_when_ArraySlice_l173_58 - _zz__zz_when_ArraySlice_l173_58_3);
      end
    end else begin
      if(when_ArraySlice_l118_58) begin
        _zz_when_ArraySlice_l173_58 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_58 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_58 = (_zz_when_ArraySlice_l118_58 <= wReg);
  assign when_ArraySlice_l173_58 = (_zz_when_ArraySlice_l173_58_1 <= _zz_when_ArraySlice_l173_58_3);
  assign when_ArraySlice_l165_59 = (_zz_when_ArraySlice_l165_59 <= selectWriteFifo);
  assign when_ArraySlice_l166_59 = (_zz_when_ArraySlice_l166_59 <= _zz_when_ArraySlice_l166_59_1);
  assign _zz_when_ArraySlice_l112_59 = (wReg % _zz__zz_when_ArraySlice_l112_59);
  assign when_ArraySlice_l112_59 = (_zz_when_ArraySlice_l112_59 != 6'h0);
  assign when_ArraySlice_l113_59 = (7'h40 <= _zz_when_ArraySlice_l113_59);
  always @(*) begin
    if(when_ArraySlice_l112_59) begin
      if(when_ArraySlice_l113_59) begin
        _zz_when_ArraySlice_l173_59 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_59 = (_zz__zz_when_ArraySlice_l173_59 - _zz__zz_when_ArraySlice_l173_59_3);
      end
    end else begin
      if(when_ArraySlice_l118_59) begin
        _zz_when_ArraySlice_l173_59 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_59 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_59 = (_zz_when_ArraySlice_l118_59 <= wReg);
  assign when_ArraySlice_l173_59 = (_zz_when_ArraySlice_l173_59_1 <= _zz_when_ArraySlice_l173_59_3);
  assign when_ArraySlice_l165_60 = (_zz_when_ArraySlice_l165_60 <= selectWriteFifo);
  assign when_ArraySlice_l166_60 = (_zz_when_ArraySlice_l166_60 <= _zz_when_ArraySlice_l166_60_1);
  assign _zz_when_ArraySlice_l112_60 = (wReg % _zz__zz_when_ArraySlice_l112_60);
  assign when_ArraySlice_l112_60 = (_zz_when_ArraySlice_l112_60 != 6'h0);
  assign when_ArraySlice_l113_60 = (7'h40 <= _zz_when_ArraySlice_l113_60);
  always @(*) begin
    if(when_ArraySlice_l112_60) begin
      if(when_ArraySlice_l113_60) begin
        _zz_when_ArraySlice_l173_60 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_60 = (_zz__zz_when_ArraySlice_l173_60 - _zz__zz_when_ArraySlice_l173_60_3);
      end
    end else begin
      if(when_ArraySlice_l118_60) begin
        _zz_when_ArraySlice_l173_60 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_60 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_60 = (_zz_when_ArraySlice_l118_60 <= wReg);
  assign when_ArraySlice_l173_60 = (_zz_when_ArraySlice_l173_60_1 <= _zz_when_ArraySlice_l173_60_3);
  assign when_ArraySlice_l165_61 = (_zz_when_ArraySlice_l165_61 <= selectWriteFifo);
  assign when_ArraySlice_l166_61 = (_zz_when_ArraySlice_l166_61 <= _zz_when_ArraySlice_l166_61_2);
  assign _zz_when_ArraySlice_l112_61 = (wReg % _zz__zz_when_ArraySlice_l112_61);
  assign when_ArraySlice_l112_61 = (_zz_when_ArraySlice_l112_61 != 6'h0);
  assign when_ArraySlice_l113_61 = (7'h40 <= _zz_when_ArraySlice_l113_61);
  always @(*) begin
    if(when_ArraySlice_l112_61) begin
      if(when_ArraySlice_l113_61) begin
        _zz_when_ArraySlice_l173_61 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_61 = (_zz__zz_when_ArraySlice_l173_61 - _zz__zz_when_ArraySlice_l173_61_3);
      end
    end else begin
      if(when_ArraySlice_l118_61) begin
        _zz_when_ArraySlice_l173_61 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_61 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_61 = (_zz_when_ArraySlice_l118_61 <= wReg);
  assign when_ArraySlice_l173_61 = (_zz_when_ArraySlice_l173_61_1 <= _zz_when_ArraySlice_l173_61_3);
  assign when_ArraySlice_l165_62 = (_zz_when_ArraySlice_l165_62 <= selectWriteFifo);
  assign when_ArraySlice_l166_62 = (_zz_when_ArraySlice_l166_62 <= _zz_when_ArraySlice_l166_62_2);
  assign _zz_when_ArraySlice_l112_62 = (wReg % _zz__zz_when_ArraySlice_l112_62);
  assign when_ArraySlice_l112_62 = (_zz_when_ArraySlice_l112_62 != 6'h0);
  assign when_ArraySlice_l113_62 = (7'h40 <= _zz_when_ArraySlice_l113_62);
  always @(*) begin
    if(when_ArraySlice_l112_62) begin
      if(when_ArraySlice_l113_62) begin
        _zz_when_ArraySlice_l173_62 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_62 = (_zz__zz_when_ArraySlice_l173_62 - _zz__zz_when_ArraySlice_l173_62_3);
      end
    end else begin
      if(when_ArraySlice_l118_62) begin
        _zz_when_ArraySlice_l173_62 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_62 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_62 = (_zz_when_ArraySlice_l118_62 <= wReg);
  assign when_ArraySlice_l173_62 = (_zz_when_ArraySlice_l173_62_1 <= _zz_when_ArraySlice_l173_62_3);
  assign when_ArraySlice_l165_63 = (_zz_when_ArraySlice_l165_63 <= selectWriteFifo);
  assign when_ArraySlice_l166_63 = (_zz_when_ArraySlice_l166_63 <= _zz_when_ArraySlice_l166_63_2);
  assign _zz_when_ArraySlice_l112_63 = (wReg % _zz__zz_when_ArraySlice_l112_63);
  assign when_ArraySlice_l112_63 = (_zz_when_ArraySlice_l112_63 != 6'h0);
  assign when_ArraySlice_l113_63 = (7'h40 <= _zz_when_ArraySlice_l113_63);
  always @(*) begin
    if(when_ArraySlice_l112_63) begin
      if(when_ArraySlice_l113_63) begin
        _zz_when_ArraySlice_l173_63 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_63 = (_zz__zz_when_ArraySlice_l173_63 - _zz__zz_when_ArraySlice_l173_63_3);
      end
    end else begin
      if(when_ArraySlice_l118_63) begin
        _zz_when_ArraySlice_l173_63 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_63 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_63 = (_zz_when_ArraySlice_l118_63 <= wReg);
  assign when_ArraySlice_l173_63 = (_zz_when_ArraySlice_l173_63_1 <= _zz_when_ArraySlice_l173_63_3);
  assign when_ArraySlice_l398_2 = (! ((((((_zz_when_ArraySlice_l398_2_1 && _zz_when_ArraySlice_l398_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l398_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l398_2_4 && _zz_when_ArraySlice_l398_2_5) && (debug_4_7 == _zz_when_ArraySlice_l398_2_6)) && (debug_5_7 == 1'b1)) && (debug_6_7 == 1'b1)) && (debug_7_7 == 1'b1))));
  assign when_ArraySlice_l401_2 = (wReg <= _zz_when_ArraySlice_l401_2_1);
  assign when_ArraySlice_l405_2 = (_zz_when_ArraySlice_l405_2_1 == 13'h0);
  assign when_ArraySlice_l409_2 = (_zz_when_ArraySlice_l409_2_1 == 7'h0);
  assign outputStreamArrayData_2_fire_2 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l410_2 = ((handshakeTimes_2_value == _zz_when_ArraySlice_l410_2_1) && outputStreamArrayData_2_fire_2);
  assign _zz_when_ArraySlice_l94_7 = (hReg % _zz__zz_when_ArraySlice_l94_7);
  assign when_ArraySlice_l94_7 = (_zz_when_ArraySlice_l94_7 != 6'h0);
  assign when_ArraySlice_l95_7 = (7'h40 <= _zz_when_ArraySlice_l95_7);
  always @(*) begin
    if(when_ArraySlice_l94_7) begin
      if(when_ArraySlice_l95_7) begin
        _zz_when_ArraySlice_l412_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_2 = (_zz__zz_when_ArraySlice_l412_2_1 - _zz__zz_when_ArraySlice_l412_2_4);
      end
    end else begin
      if(when_ArraySlice_l99_7) begin
        _zz_when_ArraySlice_l412_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_2 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_7 = (_zz_when_ArraySlice_l99_7 <= hReg);
  assign when_ArraySlice_l412_2 = (_zz_when_ArraySlice_l412_2_1 < _zz_when_ArraySlice_l412_2_4);
  always @(*) begin
    debug_0_8 = 1'b0;
    if(when_ArraySlice_l165_64) begin
      if(when_ArraySlice_l166_64) begin
        debug_0_8 = 1'b1;
      end else begin
        debug_0_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_64) begin
        debug_0_8 = 1'b1;
      end else begin
        debug_0_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_8 = 1'b0;
    if(when_ArraySlice_l165_65) begin
      if(when_ArraySlice_l166_65) begin
        debug_1_8 = 1'b1;
      end else begin
        debug_1_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_65) begin
        debug_1_8 = 1'b1;
      end else begin
        debug_1_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_8 = 1'b0;
    if(when_ArraySlice_l165_66) begin
      if(when_ArraySlice_l166_66) begin
        debug_2_8 = 1'b1;
      end else begin
        debug_2_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_66) begin
        debug_2_8 = 1'b1;
      end else begin
        debug_2_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_8 = 1'b0;
    if(when_ArraySlice_l165_67) begin
      if(when_ArraySlice_l166_67) begin
        debug_3_8 = 1'b1;
      end else begin
        debug_3_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_67) begin
        debug_3_8 = 1'b1;
      end else begin
        debug_3_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_8 = 1'b0;
    if(when_ArraySlice_l165_68) begin
      if(when_ArraySlice_l166_68) begin
        debug_4_8 = 1'b1;
      end else begin
        debug_4_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_68) begin
        debug_4_8 = 1'b1;
      end else begin
        debug_4_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_8 = 1'b0;
    if(when_ArraySlice_l165_69) begin
      if(when_ArraySlice_l166_69) begin
        debug_5_8 = 1'b1;
      end else begin
        debug_5_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_69) begin
        debug_5_8 = 1'b1;
      end else begin
        debug_5_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_8 = 1'b0;
    if(when_ArraySlice_l165_70) begin
      if(when_ArraySlice_l166_70) begin
        debug_6_8 = 1'b1;
      end else begin
        debug_6_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_70) begin
        debug_6_8 = 1'b1;
      end else begin
        debug_6_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_8 = 1'b0;
    if(when_ArraySlice_l165_71) begin
      if(when_ArraySlice_l166_71) begin
        debug_7_8 = 1'b1;
      end else begin
        debug_7_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_71) begin
        debug_7_8 = 1'b1;
      end else begin
        debug_7_8 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_64 = (_zz_when_ArraySlice_l165_64 <= selectWriteFifo);
  assign when_ArraySlice_l166_64 = (_zz_when_ArraySlice_l166_64 <= _zz_when_ArraySlice_l166_64_1);
  assign _zz_when_ArraySlice_l112_64 = (wReg % _zz__zz_when_ArraySlice_l112_64);
  assign when_ArraySlice_l112_64 = (_zz_when_ArraySlice_l112_64 != 6'h0);
  assign when_ArraySlice_l113_64 = (7'h40 <= _zz_when_ArraySlice_l113_64);
  always @(*) begin
    if(when_ArraySlice_l112_64) begin
      if(when_ArraySlice_l113_64) begin
        _zz_when_ArraySlice_l173_64 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_64 = (_zz__zz_when_ArraySlice_l173_64 - _zz__zz_when_ArraySlice_l173_64_3);
      end
    end else begin
      if(when_ArraySlice_l118_64) begin
        _zz_when_ArraySlice_l173_64 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_64 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_64 = (_zz_when_ArraySlice_l118_64 <= wReg);
  assign when_ArraySlice_l173_64 = (_zz_when_ArraySlice_l173_64_1 <= _zz_when_ArraySlice_l173_64_2);
  assign when_ArraySlice_l165_65 = (_zz_when_ArraySlice_l165_65 <= selectWriteFifo);
  assign when_ArraySlice_l166_65 = (_zz_when_ArraySlice_l166_65 <= _zz_when_ArraySlice_l166_65_1);
  assign _zz_when_ArraySlice_l112_65 = (wReg % _zz__zz_when_ArraySlice_l112_65);
  assign when_ArraySlice_l112_65 = (_zz_when_ArraySlice_l112_65 != 6'h0);
  assign when_ArraySlice_l113_65 = (7'h40 <= _zz_when_ArraySlice_l113_65);
  always @(*) begin
    if(when_ArraySlice_l112_65) begin
      if(when_ArraySlice_l113_65) begin
        _zz_when_ArraySlice_l173_65 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_65 = (_zz__zz_when_ArraySlice_l173_65 - _zz__zz_when_ArraySlice_l173_65_3);
      end
    end else begin
      if(when_ArraySlice_l118_65) begin
        _zz_when_ArraySlice_l173_65 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_65 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_65 = (_zz_when_ArraySlice_l118_65 <= wReg);
  assign when_ArraySlice_l173_65 = (_zz_when_ArraySlice_l173_65_1 <= _zz_when_ArraySlice_l173_65_3);
  assign when_ArraySlice_l165_66 = (_zz_when_ArraySlice_l165_66 <= selectWriteFifo);
  assign when_ArraySlice_l166_66 = (_zz_when_ArraySlice_l166_66 <= _zz_when_ArraySlice_l166_66_1);
  assign _zz_when_ArraySlice_l112_66 = (wReg % _zz__zz_when_ArraySlice_l112_66);
  assign when_ArraySlice_l112_66 = (_zz_when_ArraySlice_l112_66 != 6'h0);
  assign when_ArraySlice_l113_66 = (7'h40 <= _zz_when_ArraySlice_l113_66);
  always @(*) begin
    if(when_ArraySlice_l112_66) begin
      if(when_ArraySlice_l113_66) begin
        _zz_when_ArraySlice_l173_66 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_66 = (_zz__zz_when_ArraySlice_l173_66 - _zz__zz_when_ArraySlice_l173_66_3);
      end
    end else begin
      if(when_ArraySlice_l118_66) begin
        _zz_when_ArraySlice_l173_66 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_66 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_66 = (_zz_when_ArraySlice_l118_66 <= wReg);
  assign when_ArraySlice_l173_66 = (_zz_when_ArraySlice_l173_66_1 <= _zz_when_ArraySlice_l173_66_3);
  assign when_ArraySlice_l165_67 = (_zz_when_ArraySlice_l165_67 <= selectWriteFifo);
  assign when_ArraySlice_l166_67 = (_zz_when_ArraySlice_l166_67 <= _zz_when_ArraySlice_l166_67_1);
  assign _zz_when_ArraySlice_l112_67 = (wReg % _zz__zz_when_ArraySlice_l112_67);
  assign when_ArraySlice_l112_67 = (_zz_when_ArraySlice_l112_67 != 6'h0);
  assign when_ArraySlice_l113_67 = (7'h40 <= _zz_when_ArraySlice_l113_67);
  always @(*) begin
    if(when_ArraySlice_l112_67) begin
      if(when_ArraySlice_l113_67) begin
        _zz_when_ArraySlice_l173_67 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_67 = (_zz__zz_when_ArraySlice_l173_67 - _zz__zz_when_ArraySlice_l173_67_3);
      end
    end else begin
      if(when_ArraySlice_l118_67) begin
        _zz_when_ArraySlice_l173_67 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_67 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_67 = (_zz_when_ArraySlice_l118_67 <= wReg);
  assign when_ArraySlice_l173_67 = (_zz_when_ArraySlice_l173_67_1 <= _zz_when_ArraySlice_l173_67_3);
  assign when_ArraySlice_l165_68 = (_zz_when_ArraySlice_l165_68 <= selectWriteFifo);
  assign when_ArraySlice_l166_68 = (_zz_when_ArraySlice_l166_68 <= _zz_when_ArraySlice_l166_68_1);
  assign _zz_when_ArraySlice_l112_68 = (wReg % _zz__zz_when_ArraySlice_l112_68);
  assign when_ArraySlice_l112_68 = (_zz_when_ArraySlice_l112_68 != 6'h0);
  assign when_ArraySlice_l113_68 = (7'h40 <= _zz_when_ArraySlice_l113_68);
  always @(*) begin
    if(when_ArraySlice_l112_68) begin
      if(when_ArraySlice_l113_68) begin
        _zz_when_ArraySlice_l173_68 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_68 = (_zz__zz_when_ArraySlice_l173_68 - _zz__zz_when_ArraySlice_l173_68_3);
      end
    end else begin
      if(when_ArraySlice_l118_68) begin
        _zz_when_ArraySlice_l173_68 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_68 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_68 = (_zz_when_ArraySlice_l118_68 <= wReg);
  assign when_ArraySlice_l173_68 = (_zz_when_ArraySlice_l173_68_1 <= _zz_when_ArraySlice_l173_68_3);
  assign when_ArraySlice_l165_69 = (_zz_when_ArraySlice_l165_69 <= selectWriteFifo);
  assign when_ArraySlice_l166_69 = (_zz_when_ArraySlice_l166_69 <= _zz_when_ArraySlice_l166_69_2);
  assign _zz_when_ArraySlice_l112_69 = (wReg % _zz__zz_when_ArraySlice_l112_69);
  assign when_ArraySlice_l112_69 = (_zz_when_ArraySlice_l112_69 != 6'h0);
  assign when_ArraySlice_l113_69 = (7'h40 <= _zz_when_ArraySlice_l113_69);
  always @(*) begin
    if(when_ArraySlice_l112_69) begin
      if(when_ArraySlice_l113_69) begin
        _zz_when_ArraySlice_l173_69 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_69 = (_zz__zz_when_ArraySlice_l173_69 - _zz__zz_when_ArraySlice_l173_69_3);
      end
    end else begin
      if(when_ArraySlice_l118_69) begin
        _zz_when_ArraySlice_l173_69 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_69 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_69 = (_zz_when_ArraySlice_l118_69 <= wReg);
  assign when_ArraySlice_l173_69 = (_zz_when_ArraySlice_l173_69_1 <= _zz_when_ArraySlice_l173_69_3);
  assign when_ArraySlice_l165_70 = (_zz_when_ArraySlice_l165_70 <= selectWriteFifo);
  assign when_ArraySlice_l166_70 = (_zz_when_ArraySlice_l166_70 <= _zz_when_ArraySlice_l166_70_2);
  assign _zz_when_ArraySlice_l112_70 = (wReg % _zz__zz_when_ArraySlice_l112_70);
  assign when_ArraySlice_l112_70 = (_zz_when_ArraySlice_l112_70 != 6'h0);
  assign when_ArraySlice_l113_70 = (7'h40 <= _zz_when_ArraySlice_l113_70);
  always @(*) begin
    if(when_ArraySlice_l112_70) begin
      if(when_ArraySlice_l113_70) begin
        _zz_when_ArraySlice_l173_70 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_70 = (_zz__zz_when_ArraySlice_l173_70 - _zz__zz_when_ArraySlice_l173_70_3);
      end
    end else begin
      if(when_ArraySlice_l118_70) begin
        _zz_when_ArraySlice_l173_70 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_70 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_70 = (_zz_when_ArraySlice_l118_70 <= wReg);
  assign when_ArraySlice_l173_70 = (_zz_when_ArraySlice_l173_70_1 <= _zz_when_ArraySlice_l173_70_3);
  assign when_ArraySlice_l165_71 = (_zz_when_ArraySlice_l165_71 <= selectWriteFifo);
  assign when_ArraySlice_l166_71 = (_zz_when_ArraySlice_l166_71 <= _zz_when_ArraySlice_l166_71_2);
  assign _zz_when_ArraySlice_l112_71 = (wReg % _zz__zz_when_ArraySlice_l112_71);
  assign when_ArraySlice_l112_71 = (_zz_when_ArraySlice_l112_71 != 6'h0);
  assign when_ArraySlice_l113_71 = (7'h40 <= _zz_when_ArraySlice_l113_71);
  always @(*) begin
    if(when_ArraySlice_l112_71) begin
      if(when_ArraySlice_l113_71) begin
        _zz_when_ArraySlice_l173_71 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_71 = (_zz__zz_when_ArraySlice_l173_71 - _zz__zz_when_ArraySlice_l173_71_3);
      end
    end else begin
      if(when_ArraySlice_l118_71) begin
        _zz_when_ArraySlice_l173_71 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_71 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_71 = (_zz_when_ArraySlice_l118_71 <= wReg);
  assign when_ArraySlice_l173_71 = (_zz_when_ArraySlice_l173_71_1 <= _zz_when_ArraySlice_l173_71_3);
  assign when_ArraySlice_l418_2 = (! ((((((_zz_when_ArraySlice_l418_2_1 && _zz_when_ArraySlice_l418_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l418_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l418_2_4 && _zz_when_ArraySlice_l418_2_5) && (debug_4_8 == _zz_when_ArraySlice_l418_2_6)) && (debug_5_8 == 1'b1)) && (debug_6_8 == 1'b1)) && (debug_7_8 == 1'b1))));
  assign when_ArraySlice_l421_2 = (wReg <= _zz_when_ArraySlice_l421_2_1);
  assign outputStreamArrayData_2_fire_3 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l425_2 = ((_zz_when_ArraySlice_l425_2_1 == 13'h0) && outputStreamArrayData_2_fire_3);
  assign outputStreamArrayData_2_fire_4 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l436_2 = ((handshakeTimes_2_value == _zz_when_ArraySlice_l436_2_1) && outputStreamArrayData_2_fire_4);
  assign _zz_when_ArraySlice_l94_8 = (hReg % _zz__zz_when_ArraySlice_l94_8);
  assign when_ArraySlice_l94_8 = (_zz_when_ArraySlice_l94_8 != 6'h0);
  assign when_ArraySlice_l95_8 = (7'h40 <= _zz_when_ArraySlice_l95_8);
  always @(*) begin
    if(when_ArraySlice_l94_8) begin
      if(when_ArraySlice_l95_8) begin
        _zz_when_ArraySlice_l437_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_2 = (_zz__zz_when_ArraySlice_l437_2_1 - _zz__zz_when_ArraySlice_l437_2_4);
      end
    end else begin
      if(when_ArraySlice_l99_8) begin
        _zz_when_ArraySlice_l437_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_2 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_8 = (_zz_when_ArraySlice_l99_8 <= hReg);
  assign when_ArraySlice_l437_2 = (_zz_when_ArraySlice_l437_2_1 < _zz_when_ArraySlice_l437_2_4);
  always @(*) begin
    debug_0_9 = 1'b0;
    if(when_ArraySlice_l165_72) begin
      if(when_ArraySlice_l166_72) begin
        debug_0_9 = 1'b1;
      end else begin
        debug_0_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_72) begin
        debug_0_9 = 1'b1;
      end else begin
        debug_0_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_9 = 1'b0;
    if(when_ArraySlice_l165_73) begin
      if(when_ArraySlice_l166_73) begin
        debug_1_9 = 1'b1;
      end else begin
        debug_1_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_73) begin
        debug_1_9 = 1'b1;
      end else begin
        debug_1_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_9 = 1'b0;
    if(when_ArraySlice_l165_74) begin
      if(when_ArraySlice_l166_74) begin
        debug_2_9 = 1'b1;
      end else begin
        debug_2_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_74) begin
        debug_2_9 = 1'b1;
      end else begin
        debug_2_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_9 = 1'b0;
    if(when_ArraySlice_l165_75) begin
      if(when_ArraySlice_l166_75) begin
        debug_3_9 = 1'b1;
      end else begin
        debug_3_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_75) begin
        debug_3_9 = 1'b1;
      end else begin
        debug_3_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_9 = 1'b0;
    if(when_ArraySlice_l165_76) begin
      if(when_ArraySlice_l166_76) begin
        debug_4_9 = 1'b1;
      end else begin
        debug_4_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_76) begin
        debug_4_9 = 1'b1;
      end else begin
        debug_4_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_9 = 1'b0;
    if(when_ArraySlice_l165_77) begin
      if(when_ArraySlice_l166_77) begin
        debug_5_9 = 1'b1;
      end else begin
        debug_5_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_77) begin
        debug_5_9 = 1'b1;
      end else begin
        debug_5_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_9 = 1'b0;
    if(when_ArraySlice_l165_78) begin
      if(when_ArraySlice_l166_78) begin
        debug_6_9 = 1'b1;
      end else begin
        debug_6_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_78) begin
        debug_6_9 = 1'b1;
      end else begin
        debug_6_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_9 = 1'b0;
    if(when_ArraySlice_l165_79) begin
      if(when_ArraySlice_l166_79) begin
        debug_7_9 = 1'b1;
      end else begin
        debug_7_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_79) begin
        debug_7_9 = 1'b1;
      end else begin
        debug_7_9 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_72 = (_zz_when_ArraySlice_l165_72 <= selectWriteFifo);
  assign when_ArraySlice_l166_72 = (_zz_when_ArraySlice_l166_72 <= _zz_when_ArraySlice_l166_72_1);
  assign _zz_when_ArraySlice_l112_72 = (wReg % _zz__zz_when_ArraySlice_l112_72);
  assign when_ArraySlice_l112_72 = (_zz_when_ArraySlice_l112_72 != 6'h0);
  assign when_ArraySlice_l113_72 = (7'h40 <= _zz_when_ArraySlice_l113_72);
  always @(*) begin
    if(when_ArraySlice_l112_72) begin
      if(when_ArraySlice_l113_72) begin
        _zz_when_ArraySlice_l173_72 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_72 = (_zz__zz_when_ArraySlice_l173_72 - _zz__zz_when_ArraySlice_l173_72_3);
      end
    end else begin
      if(when_ArraySlice_l118_72) begin
        _zz_when_ArraySlice_l173_72 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_72 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_72 = (_zz_when_ArraySlice_l118_72 <= wReg);
  assign when_ArraySlice_l173_72 = (_zz_when_ArraySlice_l173_72_1 <= _zz_when_ArraySlice_l173_72_2);
  assign when_ArraySlice_l165_73 = (_zz_when_ArraySlice_l165_73 <= selectWriteFifo);
  assign when_ArraySlice_l166_73 = (_zz_when_ArraySlice_l166_73 <= _zz_when_ArraySlice_l166_73_1);
  assign _zz_when_ArraySlice_l112_73 = (wReg % _zz__zz_when_ArraySlice_l112_73);
  assign when_ArraySlice_l112_73 = (_zz_when_ArraySlice_l112_73 != 6'h0);
  assign when_ArraySlice_l113_73 = (7'h40 <= _zz_when_ArraySlice_l113_73);
  always @(*) begin
    if(when_ArraySlice_l112_73) begin
      if(when_ArraySlice_l113_73) begin
        _zz_when_ArraySlice_l173_73 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_73 = (_zz__zz_when_ArraySlice_l173_73 - _zz__zz_when_ArraySlice_l173_73_3);
      end
    end else begin
      if(when_ArraySlice_l118_73) begin
        _zz_when_ArraySlice_l173_73 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_73 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_73 = (_zz_when_ArraySlice_l118_73 <= wReg);
  assign when_ArraySlice_l173_73 = (_zz_when_ArraySlice_l173_73_1 <= _zz_when_ArraySlice_l173_73_3);
  assign when_ArraySlice_l165_74 = (_zz_when_ArraySlice_l165_74 <= selectWriteFifo);
  assign when_ArraySlice_l166_74 = (_zz_when_ArraySlice_l166_74 <= _zz_when_ArraySlice_l166_74_1);
  assign _zz_when_ArraySlice_l112_74 = (wReg % _zz__zz_when_ArraySlice_l112_74);
  assign when_ArraySlice_l112_74 = (_zz_when_ArraySlice_l112_74 != 6'h0);
  assign when_ArraySlice_l113_74 = (7'h40 <= _zz_when_ArraySlice_l113_74);
  always @(*) begin
    if(when_ArraySlice_l112_74) begin
      if(when_ArraySlice_l113_74) begin
        _zz_when_ArraySlice_l173_74 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_74 = (_zz__zz_when_ArraySlice_l173_74 - _zz__zz_when_ArraySlice_l173_74_3);
      end
    end else begin
      if(when_ArraySlice_l118_74) begin
        _zz_when_ArraySlice_l173_74 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_74 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_74 = (_zz_when_ArraySlice_l118_74 <= wReg);
  assign when_ArraySlice_l173_74 = (_zz_when_ArraySlice_l173_74_1 <= _zz_when_ArraySlice_l173_74_3);
  assign when_ArraySlice_l165_75 = (_zz_when_ArraySlice_l165_75 <= selectWriteFifo);
  assign when_ArraySlice_l166_75 = (_zz_when_ArraySlice_l166_75 <= _zz_when_ArraySlice_l166_75_1);
  assign _zz_when_ArraySlice_l112_75 = (wReg % _zz__zz_when_ArraySlice_l112_75);
  assign when_ArraySlice_l112_75 = (_zz_when_ArraySlice_l112_75 != 6'h0);
  assign when_ArraySlice_l113_75 = (7'h40 <= _zz_when_ArraySlice_l113_75);
  always @(*) begin
    if(when_ArraySlice_l112_75) begin
      if(when_ArraySlice_l113_75) begin
        _zz_when_ArraySlice_l173_75 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_75 = (_zz__zz_when_ArraySlice_l173_75 - _zz__zz_when_ArraySlice_l173_75_3);
      end
    end else begin
      if(when_ArraySlice_l118_75) begin
        _zz_when_ArraySlice_l173_75 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_75 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_75 = (_zz_when_ArraySlice_l118_75 <= wReg);
  assign when_ArraySlice_l173_75 = (_zz_when_ArraySlice_l173_75_1 <= _zz_when_ArraySlice_l173_75_3);
  assign when_ArraySlice_l165_76 = (_zz_when_ArraySlice_l165_76 <= selectWriteFifo);
  assign when_ArraySlice_l166_76 = (_zz_when_ArraySlice_l166_76 <= _zz_when_ArraySlice_l166_76_1);
  assign _zz_when_ArraySlice_l112_76 = (wReg % _zz__zz_when_ArraySlice_l112_76);
  assign when_ArraySlice_l112_76 = (_zz_when_ArraySlice_l112_76 != 6'h0);
  assign when_ArraySlice_l113_76 = (7'h40 <= _zz_when_ArraySlice_l113_76);
  always @(*) begin
    if(when_ArraySlice_l112_76) begin
      if(when_ArraySlice_l113_76) begin
        _zz_when_ArraySlice_l173_76 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_76 = (_zz__zz_when_ArraySlice_l173_76 - _zz__zz_when_ArraySlice_l173_76_3);
      end
    end else begin
      if(when_ArraySlice_l118_76) begin
        _zz_when_ArraySlice_l173_76 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_76 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_76 = (_zz_when_ArraySlice_l118_76 <= wReg);
  assign when_ArraySlice_l173_76 = (_zz_when_ArraySlice_l173_76_1 <= _zz_when_ArraySlice_l173_76_3);
  assign when_ArraySlice_l165_77 = (_zz_when_ArraySlice_l165_77 <= selectWriteFifo);
  assign when_ArraySlice_l166_77 = (_zz_when_ArraySlice_l166_77 <= _zz_when_ArraySlice_l166_77_2);
  assign _zz_when_ArraySlice_l112_77 = (wReg % _zz__zz_when_ArraySlice_l112_77);
  assign when_ArraySlice_l112_77 = (_zz_when_ArraySlice_l112_77 != 6'h0);
  assign when_ArraySlice_l113_77 = (7'h40 <= _zz_when_ArraySlice_l113_77);
  always @(*) begin
    if(when_ArraySlice_l112_77) begin
      if(when_ArraySlice_l113_77) begin
        _zz_when_ArraySlice_l173_77 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_77 = (_zz__zz_when_ArraySlice_l173_77 - _zz__zz_when_ArraySlice_l173_77_3);
      end
    end else begin
      if(when_ArraySlice_l118_77) begin
        _zz_when_ArraySlice_l173_77 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_77 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_77 = (_zz_when_ArraySlice_l118_77 <= wReg);
  assign when_ArraySlice_l173_77 = (_zz_when_ArraySlice_l173_77_1 <= _zz_when_ArraySlice_l173_77_3);
  assign when_ArraySlice_l165_78 = (_zz_when_ArraySlice_l165_78 <= selectWriteFifo);
  assign when_ArraySlice_l166_78 = (_zz_when_ArraySlice_l166_78 <= _zz_when_ArraySlice_l166_78_2);
  assign _zz_when_ArraySlice_l112_78 = (wReg % _zz__zz_when_ArraySlice_l112_78);
  assign when_ArraySlice_l112_78 = (_zz_when_ArraySlice_l112_78 != 6'h0);
  assign when_ArraySlice_l113_78 = (7'h40 <= _zz_when_ArraySlice_l113_78);
  always @(*) begin
    if(when_ArraySlice_l112_78) begin
      if(when_ArraySlice_l113_78) begin
        _zz_when_ArraySlice_l173_78 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_78 = (_zz__zz_when_ArraySlice_l173_78 - _zz__zz_when_ArraySlice_l173_78_3);
      end
    end else begin
      if(when_ArraySlice_l118_78) begin
        _zz_when_ArraySlice_l173_78 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_78 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_78 = (_zz_when_ArraySlice_l118_78 <= wReg);
  assign when_ArraySlice_l173_78 = (_zz_when_ArraySlice_l173_78_1 <= _zz_when_ArraySlice_l173_78_3);
  assign when_ArraySlice_l165_79 = (_zz_when_ArraySlice_l165_79 <= selectWriteFifo);
  assign when_ArraySlice_l166_79 = (_zz_when_ArraySlice_l166_79 <= _zz_when_ArraySlice_l166_79_2);
  assign _zz_when_ArraySlice_l112_79 = (wReg % _zz__zz_when_ArraySlice_l112_79);
  assign when_ArraySlice_l112_79 = (_zz_when_ArraySlice_l112_79 != 6'h0);
  assign when_ArraySlice_l113_79 = (7'h40 <= _zz_when_ArraySlice_l113_79);
  always @(*) begin
    if(when_ArraySlice_l112_79) begin
      if(when_ArraySlice_l113_79) begin
        _zz_when_ArraySlice_l173_79 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_79 = (_zz__zz_when_ArraySlice_l173_79 - _zz__zz_when_ArraySlice_l173_79_3);
      end
    end else begin
      if(when_ArraySlice_l118_79) begin
        _zz_when_ArraySlice_l173_79 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_79 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_79 = (_zz_when_ArraySlice_l118_79 <= wReg);
  assign when_ArraySlice_l173_79 = (_zz_when_ArraySlice_l173_79_1 <= _zz_when_ArraySlice_l173_79_3);
  assign when_ArraySlice_l444_2 = (! ((((((_zz_when_ArraySlice_l444_2_1 && _zz_when_ArraySlice_l444_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l444_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l444_2_4 && _zz_when_ArraySlice_l444_2_5) && (debug_4_9 == _zz_when_ArraySlice_l444_2_6)) && (debug_5_9 == 1'b1)) && (debug_6_9 == 1'b1)) && (debug_7_9 == 1'b1))));
  assign outputStreamArrayData_2_fire_5 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l448_2 = ((_zz_when_ArraySlice_l448_2_1 == 13'h0) && outputStreamArrayData_2_fire_5);
  assign when_ArraySlice_l434_2 = (allowPadding_2 && (wReg <= _zz_when_ArraySlice_l434_2_1));
  assign outputStreamArrayData_2_fire_6 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l455_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l455_2_1);
  assign when_ArraySlice_l373_3 = (_zz_when_ArraySlice_l373_3 < wReg);
  assign when_ArraySlice_l374_3 = ((! holdReadOp_3) && (_zz_when_ArraySlice_l374_3_1 != 7'h0));
  assign _zz_outputStreamArrayData_3_valid = (selectReadFifo_3 + _zz__zz_outputStreamArrayData_3_valid);
  assign _zz_6 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_3_valid);
  assign _zz_io_pop_ready_3 = outputStreamArrayData_3_ready;
  assign when_ArraySlice_l379_3 = (! holdReadOp_3);
  assign outputStreamArrayData_3_fire = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l380_3 = ((_zz_when_ArraySlice_l380_3_1 < _zz_when_ArraySlice_l380_3_3) && outputStreamArrayData_3_fire);
  assign when_ArraySlice_l381_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l381_3_1);
  assign when_ArraySlice_l384_3 = (_zz_when_ArraySlice_l384_3_1 == 13'h0);
  assign outputStreamArrayData_3_fire_1 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l389_3 = ((_zz_when_ArraySlice_l389_3_1 == _zz_when_ArraySlice_l389_3_5) && outputStreamArrayData_3_fire_1);
  assign when_ArraySlice_l390_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l390_3_1);
  assign _zz_when_ArraySlice_l94_9 = (hReg % _zz__zz_when_ArraySlice_l94_9);
  assign when_ArraySlice_l94_9 = (_zz_when_ArraySlice_l94_9 != 6'h0);
  assign when_ArraySlice_l95_9 = (7'h40 <= _zz_when_ArraySlice_l95_9);
  always @(*) begin
    if(when_ArraySlice_l94_9) begin
      if(when_ArraySlice_l95_9) begin
        _zz_when_ArraySlice_l392_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_3 = (_zz__zz_when_ArraySlice_l392_3_1 - _zz__zz_when_ArraySlice_l392_3_4);
      end
    end else begin
      if(when_ArraySlice_l99_9) begin
        _zz_when_ArraySlice_l392_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_3 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_9 = (_zz_when_ArraySlice_l99_9 <= hReg);
  assign when_ArraySlice_l392_3 = (_zz_when_ArraySlice_l392_3_1 < _zz_when_ArraySlice_l392_3_4);
  always @(*) begin
    debug_0_10 = 1'b0;
    if(when_ArraySlice_l165_80) begin
      if(when_ArraySlice_l166_80) begin
        debug_0_10 = 1'b1;
      end else begin
        debug_0_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_80) begin
        debug_0_10 = 1'b1;
      end else begin
        debug_0_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_10 = 1'b0;
    if(when_ArraySlice_l165_81) begin
      if(when_ArraySlice_l166_81) begin
        debug_1_10 = 1'b1;
      end else begin
        debug_1_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_81) begin
        debug_1_10 = 1'b1;
      end else begin
        debug_1_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_10 = 1'b0;
    if(when_ArraySlice_l165_82) begin
      if(when_ArraySlice_l166_82) begin
        debug_2_10 = 1'b1;
      end else begin
        debug_2_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_82) begin
        debug_2_10 = 1'b1;
      end else begin
        debug_2_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_10 = 1'b0;
    if(when_ArraySlice_l165_83) begin
      if(when_ArraySlice_l166_83) begin
        debug_3_10 = 1'b1;
      end else begin
        debug_3_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_83) begin
        debug_3_10 = 1'b1;
      end else begin
        debug_3_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_10 = 1'b0;
    if(when_ArraySlice_l165_84) begin
      if(when_ArraySlice_l166_84) begin
        debug_4_10 = 1'b1;
      end else begin
        debug_4_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_84) begin
        debug_4_10 = 1'b1;
      end else begin
        debug_4_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_10 = 1'b0;
    if(when_ArraySlice_l165_85) begin
      if(when_ArraySlice_l166_85) begin
        debug_5_10 = 1'b1;
      end else begin
        debug_5_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_85) begin
        debug_5_10 = 1'b1;
      end else begin
        debug_5_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_10 = 1'b0;
    if(when_ArraySlice_l165_86) begin
      if(when_ArraySlice_l166_86) begin
        debug_6_10 = 1'b1;
      end else begin
        debug_6_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_86) begin
        debug_6_10 = 1'b1;
      end else begin
        debug_6_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_10 = 1'b0;
    if(when_ArraySlice_l165_87) begin
      if(when_ArraySlice_l166_87) begin
        debug_7_10 = 1'b1;
      end else begin
        debug_7_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_87) begin
        debug_7_10 = 1'b1;
      end else begin
        debug_7_10 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_80 = (_zz_when_ArraySlice_l165_80 <= selectWriteFifo);
  assign when_ArraySlice_l166_80 = (_zz_when_ArraySlice_l166_80 <= _zz_when_ArraySlice_l166_80_1);
  assign _zz_when_ArraySlice_l112_80 = (wReg % _zz__zz_when_ArraySlice_l112_80);
  assign when_ArraySlice_l112_80 = (_zz_when_ArraySlice_l112_80 != 6'h0);
  assign when_ArraySlice_l113_80 = (7'h40 <= _zz_when_ArraySlice_l113_80);
  always @(*) begin
    if(when_ArraySlice_l112_80) begin
      if(when_ArraySlice_l113_80) begin
        _zz_when_ArraySlice_l173_80 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_80 = (_zz__zz_when_ArraySlice_l173_80 - _zz__zz_when_ArraySlice_l173_80_3);
      end
    end else begin
      if(when_ArraySlice_l118_80) begin
        _zz_when_ArraySlice_l173_80 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_80 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_80 = (_zz_when_ArraySlice_l118_80 <= wReg);
  assign when_ArraySlice_l173_80 = (_zz_when_ArraySlice_l173_80_1 <= _zz_when_ArraySlice_l173_80_2);
  assign when_ArraySlice_l165_81 = (_zz_when_ArraySlice_l165_81 <= selectWriteFifo);
  assign when_ArraySlice_l166_81 = (_zz_when_ArraySlice_l166_81 <= _zz_when_ArraySlice_l166_81_1);
  assign _zz_when_ArraySlice_l112_81 = (wReg % _zz__zz_when_ArraySlice_l112_81);
  assign when_ArraySlice_l112_81 = (_zz_when_ArraySlice_l112_81 != 6'h0);
  assign when_ArraySlice_l113_81 = (7'h40 <= _zz_when_ArraySlice_l113_81);
  always @(*) begin
    if(when_ArraySlice_l112_81) begin
      if(when_ArraySlice_l113_81) begin
        _zz_when_ArraySlice_l173_81 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_81 = (_zz__zz_when_ArraySlice_l173_81 - _zz__zz_when_ArraySlice_l173_81_3);
      end
    end else begin
      if(when_ArraySlice_l118_81) begin
        _zz_when_ArraySlice_l173_81 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_81 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_81 = (_zz_when_ArraySlice_l118_81 <= wReg);
  assign when_ArraySlice_l173_81 = (_zz_when_ArraySlice_l173_81_1 <= _zz_when_ArraySlice_l173_81_3);
  assign when_ArraySlice_l165_82 = (_zz_when_ArraySlice_l165_82 <= selectWriteFifo);
  assign when_ArraySlice_l166_82 = (_zz_when_ArraySlice_l166_82 <= _zz_when_ArraySlice_l166_82_1);
  assign _zz_when_ArraySlice_l112_82 = (wReg % _zz__zz_when_ArraySlice_l112_82);
  assign when_ArraySlice_l112_82 = (_zz_when_ArraySlice_l112_82 != 6'h0);
  assign when_ArraySlice_l113_82 = (7'h40 <= _zz_when_ArraySlice_l113_82);
  always @(*) begin
    if(when_ArraySlice_l112_82) begin
      if(when_ArraySlice_l113_82) begin
        _zz_when_ArraySlice_l173_82 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_82 = (_zz__zz_when_ArraySlice_l173_82 - _zz__zz_when_ArraySlice_l173_82_3);
      end
    end else begin
      if(when_ArraySlice_l118_82) begin
        _zz_when_ArraySlice_l173_82 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_82 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_82 = (_zz_when_ArraySlice_l118_82 <= wReg);
  assign when_ArraySlice_l173_82 = (_zz_when_ArraySlice_l173_82_1 <= _zz_when_ArraySlice_l173_82_3);
  assign when_ArraySlice_l165_83 = (_zz_when_ArraySlice_l165_83 <= selectWriteFifo);
  assign when_ArraySlice_l166_83 = (_zz_when_ArraySlice_l166_83 <= _zz_when_ArraySlice_l166_83_1);
  assign _zz_when_ArraySlice_l112_83 = (wReg % _zz__zz_when_ArraySlice_l112_83);
  assign when_ArraySlice_l112_83 = (_zz_when_ArraySlice_l112_83 != 6'h0);
  assign when_ArraySlice_l113_83 = (7'h40 <= _zz_when_ArraySlice_l113_83);
  always @(*) begin
    if(when_ArraySlice_l112_83) begin
      if(when_ArraySlice_l113_83) begin
        _zz_when_ArraySlice_l173_83 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_83 = (_zz__zz_when_ArraySlice_l173_83 - _zz__zz_when_ArraySlice_l173_83_3);
      end
    end else begin
      if(when_ArraySlice_l118_83) begin
        _zz_when_ArraySlice_l173_83 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_83 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_83 = (_zz_when_ArraySlice_l118_83 <= wReg);
  assign when_ArraySlice_l173_83 = (_zz_when_ArraySlice_l173_83_1 <= _zz_when_ArraySlice_l173_83_3);
  assign when_ArraySlice_l165_84 = (_zz_when_ArraySlice_l165_84 <= selectWriteFifo);
  assign when_ArraySlice_l166_84 = (_zz_when_ArraySlice_l166_84 <= _zz_when_ArraySlice_l166_84_1);
  assign _zz_when_ArraySlice_l112_84 = (wReg % _zz__zz_when_ArraySlice_l112_84);
  assign when_ArraySlice_l112_84 = (_zz_when_ArraySlice_l112_84 != 6'h0);
  assign when_ArraySlice_l113_84 = (7'h40 <= _zz_when_ArraySlice_l113_84);
  always @(*) begin
    if(when_ArraySlice_l112_84) begin
      if(when_ArraySlice_l113_84) begin
        _zz_when_ArraySlice_l173_84 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_84 = (_zz__zz_when_ArraySlice_l173_84 - _zz__zz_when_ArraySlice_l173_84_3);
      end
    end else begin
      if(when_ArraySlice_l118_84) begin
        _zz_when_ArraySlice_l173_84 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_84 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_84 = (_zz_when_ArraySlice_l118_84 <= wReg);
  assign when_ArraySlice_l173_84 = (_zz_when_ArraySlice_l173_84_1 <= _zz_when_ArraySlice_l173_84_3);
  assign when_ArraySlice_l165_85 = (_zz_when_ArraySlice_l165_85 <= selectWriteFifo);
  assign when_ArraySlice_l166_85 = (_zz_when_ArraySlice_l166_85 <= _zz_when_ArraySlice_l166_85_2);
  assign _zz_when_ArraySlice_l112_85 = (wReg % _zz__zz_when_ArraySlice_l112_85);
  assign when_ArraySlice_l112_85 = (_zz_when_ArraySlice_l112_85 != 6'h0);
  assign when_ArraySlice_l113_85 = (7'h40 <= _zz_when_ArraySlice_l113_85);
  always @(*) begin
    if(when_ArraySlice_l112_85) begin
      if(when_ArraySlice_l113_85) begin
        _zz_when_ArraySlice_l173_85 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_85 = (_zz__zz_when_ArraySlice_l173_85 - _zz__zz_when_ArraySlice_l173_85_3);
      end
    end else begin
      if(when_ArraySlice_l118_85) begin
        _zz_when_ArraySlice_l173_85 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_85 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_85 = (_zz_when_ArraySlice_l118_85 <= wReg);
  assign when_ArraySlice_l173_85 = (_zz_when_ArraySlice_l173_85_1 <= _zz_when_ArraySlice_l173_85_3);
  assign when_ArraySlice_l165_86 = (_zz_when_ArraySlice_l165_86 <= selectWriteFifo);
  assign when_ArraySlice_l166_86 = (_zz_when_ArraySlice_l166_86 <= _zz_when_ArraySlice_l166_86_2);
  assign _zz_when_ArraySlice_l112_86 = (wReg % _zz__zz_when_ArraySlice_l112_86);
  assign when_ArraySlice_l112_86 = (_zz_when_ArraySlice_l112_86 != 6'h0);
  assign when_ArraySlice_l113_86 = (7'h40 <= _zz_when_ArraySlice_l113_86);
  always @(*) begin
    if(when_ArraySlice_l112_86) begin
      if(when_ArraySlice_l113_86) begin
        _zz_when_ArraySlice_l173_86 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_86 = (_zz__zz_when_ArraySlice_l173_86 - _zz__zz_when_ArraySlice_l173_86_3);
      end
    end else begin
      if(when_ArraySlice_l118_86) begin
        _zz_when_ArraySlice_l173_86 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_86 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_86 = (_zz_when_ArraySlice_l118_86 <= wReg);
  assign when_ArraySlice_l173_86 = (_zz_when_ArraySlice_l173_86_1 <= _zz_when_ArraySlice_l173_86_3);
  assign when_ArraySlice_l165_87 = (_zz_when_ArraySlice_l165_87 <= selectWriteFifo);
  assign when_ArraySlice_l166_87 = (_zz_when_ArraySlice_l166_87 <= _zz_when_ArraySlice_l166_87_2);
  assign _zz_when_ArraySlice_l112_87 = (wReg % _zz__zz_when_ArraySlice_l112_87);
  assign when_ArraySlice_l112_87 = (_zz_when_ArraySlice_l112_87 != 6'h0);
  assign when_ArraySlice_l113_87 = (7'h40 <= _zz_when_ArraySlice_l113_87);
  always @(*) begin
    if(when_ArraySlice_l112_87) begin
      if(when_ArraySlice_l113_87) begin
        _zz_when_ArraySlice_l173_87 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_87 = (_zz__zz_when_ArraySlice_l173_87 - _zz__zz_when_ArraySlice_l173_87_3);
      end
    end else begin
      if(when_ArraySlice_l118_87) begin
        _zz_when_ArraySlice_l173_87 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_87 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_87 = (_zz_when_ArraySlice_l118_87 <= wReg);
  assign when_ArraySlice_l173_87 = (_zz_when_ArraySlice_l173_87_1 <= _zz_when_ArraySlice_l173_87_3);
  assign when_ArraySlice_l398_3 = (! ((((((_zz_when_ArraySlice_l398_3_1 && _zz_when_ArraySlice_l398_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l398_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l398_3_4 && _zz_when_ArraySlice_l398_3_5) && (debug_4_10 == _zz_when_ArraySlice_l398_3_6)) && (debug_5_10 == 1'b1)) && (debug_6_10 == 1'b1)) && (debug_7_10 == 1'b1))));
  assign when_ArraySlice_l401_3 = (wReg <= _zz_when_ArraySlice_l401_3_1);
  assign when_ArraySlice_l405_3 = (_zz_when_ArraySlice_l405_3_1 == 13'h0);
  assign when_ArraySlice_l409_3 = (_zz_when_ArraySlice_l409_3_1 == 7'h0);
  assign outputStreamArrayData_3_fire_2 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l410_3 = ((handshakeTimes_3_value == _zz_when_ArraySlice_l410_3_1) && outputStreamArrayData_3_fire_2);
  assign _zz_when_ArraySlice_l94_10 = (hReg % _zz__zz_when_ArraySlice_l94_10);
  assign when_ArraySlice_l94_10 = (_zz_when_ArraySlice_l94_10 != 6'h0);
  assign when_ArraySlice_l95_10 = (7'h40 <= _zz_when_ArraySlice_l95_10);
  always @(*) begin
    if(when_ArraySlice_l94_10) begin
      if(when_ArraySlice_l95_10) begin
        _zz_when_ArraySlice_l412_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_3 = (_zz__zz_when_ArraySlice_l412_3_1 - _zz__zz_when_ArraySlice_l412_3_4);
      end
    end else begin
      if(when_ArraySlice_l99_10) begin
        _zz_when_ArraySlice_l412_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_3 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_10 = (_zz_when_ArraySlice_l99_10 <= hReg);
  assign when_ArraySlice_l412_3 = (_zz_when_ArraySlice_l412_3_1 < _zz_when_ArraySlice_l412_3_4);
  always @(*) begin
    debug_0_11 = 1'b0;
    if(when_ArraySlice_l165_88) begin
      if(when_ArraySlice_l166_88) begin
        debug_0_11 = 1'b1;
      end else begin
        debug_0_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_88) begin
        debug_0_11 = 1'b1;
      end else begin
        debug_0_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_11 = 1'b0;
    if(when_ArraySlice_l165_89) begin
      if(when_ArraySlice_l166_89) begin
        debug_1_11 = 1'b1;
      end else begin
        debug_1_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_89) begin
        debug_1_11 = 1'b1;
      end else begin
        debug_1_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_11 = 1'b0;
    if(when_ArraySlice_l165_90) begin
      if(when_ArraySlice_l166_90) begin
        debug_2_11 = 1'b1;
      end else begin
        debug_2_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_90) begin
        debug_2_11 = 1'b1;
      end else begin
        debug_2_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_11 = 1'b0;
    if(when_ArraySlice_l165_91) begin
      if(when_ArraySlice_l166_91) begin
        debug_3_11 = 1'b1;
      end else begin
        debug_3_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_91) begin
        debug_3_11 = 1'b1;
      end else begin
        debug_3_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_11 = 1'b0;
    if(when_ArraySlice_l165_92) begin
      if(when_ArraySlice_l166_92) begin
        debug_4_11 = 1'b1;
      end else begin
        debug_4_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_92) begin
        debug_4_11 = 1'b1;
      end else begin
        debug_4_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_11 = 1'b0;
    if(when_ArraySlice_l165_93) begin
      if(when_ArraySlice_l166_93) begin
        debug_5_11 = 1'b1;
      end else begin
        debug_5_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_93) begin
        debug_5_11 = 1'b1;
      end else begin
        debug_5_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_11 = 1'b0;
    if(when_ArraySlice_l165_94) begin
      if(when_ArraySlice_l166_94) begin
        debug_6_11 = 1'b1;
      end else begin
        debug_6_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_94) begin
        debug_6_11 = 1'b1;
      end else begin
        debug_6_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_11 = 1'b0;
    if(when_ArraySlice_l165_95) begin
      if(when_ArraySlice_l166_95) begin
        debug_7_11 = 1'b1;
      end else begin
        debug_7_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_95) begin
        debug_7_11 = 1'b1;
      end else begin
        debug_7_11 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_88 = (_zz_when_ArraySlice_l165_88 <= selectWriteFifo);
  assign when_ArraySlice_l166_88 = (_zz_when_ArraySlice_l166_88 <= _zz_when_ArraySlice_l166_88_1);
  assign _zz_when_ArraySlice_l112_88 = (wReg % _zz__zz_when_ArraySlice_l112_88);
  assign when_ArraySlice_l112_88 = (_zz_when_ArraySlice_l112_88 != 6'h0);
  assign when_ArraySlice_l113_88 = (7'h40 <= _zz_when_ArraySlice_l113_88);
  always @(*) begin
    if(when_ArraySlice_l112_88) begin
      if(when_ArraySlice_l113_88) begin
        _zz_when_ArraySlice_l173_88 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_88 = (_zz__zz_when_ArraySlice_l173_88 - _zz__zz_when_ArraySlice_l173_88_3);
      end
    end else begin
      if(when_ArraySlice_l118_88) begin
        _zz_when_ArraySlice_l173_88 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_88 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_88 = (_zz_when_ArraySlice_l118_88 <= wReg);
  assign when_ArraySlice_l173_88 = (_zz_when_ArraySlice_l173_88_1 <= _zz_when_ArraySlice_l173_88_2);
  assign when_ArraySlice_l165_89 = (_zz_when_ArraySlice_l165_89 <= selectWriteFifo);
  assign when_ArraySlice_l166_89 = (_zz_when_ArraySlice_l166_89 <= _zz_when_ArraySlice_l166_89_1);
  assign _zz_when_ArraySlice_l112_89 = (wReg % _zz__zz_when_ArraySlice_l112_89);
  assign when_ArraySlice_l112_89 = (_zz_when_ArraySlice_l112_89 != 6'h0);
  assign when_ArraySlice_l113_89 = (7'h40 <= _zz_when_ArraySlice_l113_89);
  always @(*) begin
    if(when_ArraySlice_l112_89) begin
      if(when_ArraySlice_l113_89) begin
        _zz_when_ArraySlice_l173_89 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_89 = (_zz__zz_when_ArraySlice_l173_89 - _zz__zz_when_ArraySlice_l173_89_3);
      end
    end else begin
      if(when_ArraySlice_l118_89) begin
        _zz_when_ArraySlice_l173_89 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_89 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_89 = (_zz_when_ArraySlice_l118_89 <= wReg);
  assign when_ArraySlice_l173_89 = (_zz_when_ArraySlice_l173_89_1 <= _zz_when_ArraySlice_l173_89_3);
  assign when_ArraySlice_l165_90 = (_zz_when_ArraySlice_l165_90 <= selectWriteFifo);
  assign when_ArraySlice_l166_90 = (_zz_when_ArraySlice_l166_90 <= _zz_when_ArraySlice_l166_90_1);
  assign _zz_when_ArraySlice_l112_90 = (wReg % _zz__zz_when_ArraySlice_l112_90);
  assign when_ArraySlice_l112_90 = (_zz_when_ArraySlice_l112_90 != 6'h0);
  assign when_ArraySlice_l113_90 = (7'h40 <= _zz_when_ArraySlice_l113_90);
  always @(*) begin
    if(when_ArraySlice_l112_90) begin
      if(when_ArraySlice_l113_90) begin
        _zz_when_ArraySlice_l173_90 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_90 = (_zz__zz_when_ArraySlice_l173_90 - _zz__zz_when_ArraySlice_l173_90_3);
      end
    end else begin
      if(when_ArraySlice_l118_90) begin
        _zz_when_ArraySlice_l173_90 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_90 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_90 = (_zz_when_ArraySlice_l118_90 <= wReg);
  assign when_ArraySlice_l173_90 = (_zz_when_ArraySlice_l173_90_1 <= _zz_when_ArraySlice_l173_90_3);
  assign when_ArraySlice_l165_91 = (_zz_when_ArraySlice_l165_91 <= selectWriteFifo);
  assign when_ArraySlice_l166_91 = (_zz_when_ArraySlice_l166_91 <= _zz_when_ArraySlice_l166_91_1);
  assign _zz_when_ArraySlice_l112_91 = (wReg % _zz__zz_when_ArraySlice_l112_91);
  assign when_ArraySlice_l112_91 = (_zz_when_ArraySlice_l112_91 != 6'h0);
  assign when_ArraySlice_l113_91 = (7'h40 <= _zz_when_ArraySlice_l113_91);
  always @(*) begin
    if(when_ArraySlice_l112_91) begin
      if(when_ArraySlice_l113_91) begin
        _zz_when_ArraySlice_l173_91 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_91 = (_zz__zz_when_ArraySlice_l173_91 - _zz__zz_when_ArraySlice_l173_91_3);
      end
    end else begin
      if(when_ArraySlice_l118_91) begin
        _zz_when_ArraySlice_l173_91 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_91 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_91 = (_zz_when_ArraySlice_l118_91 <= wReg);
  assign when_ArraySlice_l173_91 = (_zz_when_ArraySlice_l173_91_1 <= _zz_when_ArraySlice_l173_91_3);
  assign when_ArraySlice_l165_92 = (_zz_when_ArraySlice_l165_92 <= selectWriteFifo);
  assign when_ArraySlice_l166_92 = (_zz_when_ArraySlice_l166_92 <= _zz_when_ArraySlice_l166_92_1);
  assign _zz_when_ArraySlice_l112_92 = (wReg % _zz__zz_when_ArraySlice_l112_92);
  assign when_ArraySlice_l112_92 = (_zz_when_ArraySlice_l112_92 != 6'h0);
  assign when_ArraySlice_l113_92 = (7'h40 <= _zz_when_ArraySlice_l113_92);
  always @(*) begin
    if(when_ArraySlice_l112_92) begin
      if(when_ArraySlice_l113_92) begin
        _zz_when_ArraySlice_l173_92 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_92 = (_zz__zz_when_ArraySlice_l173_92 - _zz__zz_when_ArraySlice_l173_92_3);
      end
    end else begin
      if(when_ArraySlice_l118_92) begin
        _zz_when_ArraySlice_l173_92 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_92 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_92 = (_zz_when_ArraySlice_l118_92 <= wReg);
  assign when_ArraySlice_l173_92 = (_zz_when_ArraySlice_l173_92_1 <= _zz_when_ArraySlice_l173_92_3);
  assign when_ArraySlice_l165_93 = (_zz_when_ArraySlice_l165_93 <= selectWriteFifo);
  assign when_ArraySlice_l166_93 = (_zz_when_ArraySlice_l166_93 <= _zz_when_ArraySlice_l166_93_2);
  assign _zz_when_ArraySlice_l112_93 = (wReg % _zz__zz_when_ArraySlice_l112_93);
  assign when_ArraySlice_l112_93 = (_zz_when_ArraySlice_l112_93 != 6'h0);
  assign when_ArraySlice_l113_93 = (7'h40 <= _zz_when_ArraySlice_l113_93);
  always @(*) begin
    if(when_ArraySlice_l112_93) begin
      if(when_ArraySlice_l113_93) begin
        _zz_when_ArraySlice_l173_93 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_93 = (_zz__zz_when_ArraySlice_l173_93 - _zz__zz_when_ArraySlice_l173_93_3);
      end
    end else begin
      if(when_ArraySlice_l118_93) begin
        _zz_when_ArraySlice_l173_93 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_93 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_93 = (_zz_when_ArraySlice_l118_93 <= wReg);
  assign when_ArraySlice_l173_93 = (_zz_when_ArraySlice_l173_93_1 <= _zz_when_ArraySlice_l173_93_3);
  assign when_ArraySlice_l165_94 = (_zz_when_ArraySlice_l165_94 <= selectWriteFifo);
  assign when_ArraySlice_l166_94 = (_zz_when_ArraySlice_l166_94 <= _zz_when_ArraySlice_l166_94_2);
  assign _zz_when_ArraySlice_l112_94 = (wReg % _zz__zz_when_ArraySlice_l112_94);
  assign when_ArraySlice_l112_94 = (_zz_when_ArraySlice_l112_94 != 6'h0);
  assign when_ArraySlice_l113_94 = (7'h40 <= _zz_when_ArraySlice_l113_94);
  always @(*) begin
    if(when_ArraySlice_l112_94) begin
      if(when_ArraySlice_l113_94) begin
        _zz_when_ArraySlice_l173_94 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_94 = (_zz__zz_when_ArraySlice_l173_94 - _zz__zz_when_ArraySlice_l173_94_3);
      end
    end else begin
      if(when_ArraySlice_l118_94) begin
        _zz_when_ArraySlice_l173_94 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_94 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_94 = (_zz_when_ArraySlice_l118_94 <= wReg);
  assign when_ArraySlice_l173_94 = (_zz_when_ArraySlice_l173_94_1 <= _zz_when_ArraySlice_l173_94_3);
  assign when_ArraySlice_l165_95 = (_zz_when_ArraySlice_l165_95 <= selectWriteFifo);
  assign when_ArraySlice_l166_95 = (_zz_when_ArraySlice_l166_95 <= _zz_when_ArraySlice_l166_95_2);
  assign _zz_when_ArraySlice_l112_95 = (wReg % _zz__zz_when_ArraySlice_l112_95);
  assign when_ArraySlice_l112_95 = (_zz_when_ArraySlice_l112_95 != 6'h0);
  assign when_ArraySlice_l113_95 = (7'h40 <= _zz_when_ArraySlice_l113_95);
  always @(*) begin
    if(when_ArraySlice_l112_95) begin
      if(when_ArraySlice_l113_95) begin
        _zz_when_ArraySlice_l173_95 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_95 = (_zz__zz_when_ArraySlice_l173_95 - _zz__zz_when_ArraySlice_l173_95_3);
      end
    end else begin
      if(when_ArraySlice_l118_95) begin
        _zz_when_ArraySlice_l173_95 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_95 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_95 = (_zz_when_ArraySlice_l118_95 <= wReg);
  assign when_ArraySlice_l173_95 = (_zz_when_ArraySlice_l173_95_1 <= _zz_when_ArraySlice_l173_95_3);
  assign when_ArraySlice_l418_3 = (! ((((((_zz_when_ArraySlice_l418_3_1 && _zz_when_ArraySlice_l418_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l418_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l418_3_4 && _zz_when_ArraySlice_l418_3_5) && (debug_4_11 == _zz_when_ArraySlice_l418_3_6)) && (debug_5_11 == 1'b1)) && (debug_6_11 == 1'b1)) && (debug_7_11 == 1'b1))));
  assign when_ArraySlice_l421_3 = (wReg <= _zz_when_ArraySlice_l421_3_1);
  assign outputStreamArrayData_3_fire_3 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l425_3 = ((_zz_when_ArraySlice_l425_3_1 == 13'h0) && outputStreamArrayData_3_fire_3);
  assign outputStreamArrayData_3_fire_4 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l436_3 = ((handshakeTimes_3_value == _zz_when_ArraySlice_l436_3_1) && outputStreamArrayData_3_fire_4);
  assign _zz_when_ArraySlice_l94_11 = (hReg % _zz__zz_when_ArraySlice_l94_11);
  assign when_ArraySlice_l94_11 = (_zz_when_ArraySlice_l94_11 != 6'h0);
  assign when_ArraySlice_l95_11 = (7'h40 <= _zz_when_ArraySlice_l95_11);
  always @(*) begin
    if(when_ArraySlice_l94_11) begin
      if(when_ArraySlice_l95_11) begin
        _zz_when_ArraySlice_l437_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_3 = (_zz__zz_when_ArraySlice_l437_3_1 - _zz__zz_when_ArraySlice_l437_3_4);
      end
    end else begin
      if(when_ArraySlice_l99_11) begin
        _zz_when_ArraySlice_l437_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_3 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_11 = (_zz_when_ArraySlice_l99_11 <= hReg);
  assign when_ArraySlice_l437_3 = (_zz_when_ArraySlice_l437_3_1 < _zz_when_ArraySlice_l437_3_4);
  always @(*) begin
    debug_0_12 = 1'b0;
    if(when_ArraySlice_l165_96) begin
      if(when_ArraySlice_l166_96) begin
        debug_0_12 = 1'b1;
      end else begin
        debug_0_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_96) begin
        debug_0_12 = 1'b1;
      end else begin
        debug_0_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_12 = 1'b0;
    if(when_ArraySlice_l165_97) begin
      if(when_ArraySlice_l166_97) begin
        debug_1_12 = 1'b1;
      end else begin
        debug_1_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_97) begin
        debug_1_12 = 1'b1;
      end else begin
        debug_1_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_12 = 1'b0;
    if(when_ArraySlice_l165_98) begin
      if(when_ArraySlice_l166_98) begin
        debug_2_12 = 1'b1;
      end else begin
        debug_2_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_98) begin
        debug_2_12 = 1'b1;
      end else begin
        debug_2_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_12 = 1'b0;
    if(when_ArraySlice_l165_99) begin
      if(when_ArraySlice_l166_99) begin
        debug_3_12 = 1'b1;
      end else begin
        debug_3_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_99) begin
        debug_3_12 = 1'b1;
      end else begin
        debug_3_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_12 = 1'b0;
    if(when_ArraySlice_l165_100) begin
      if(when_ArraySlice_l166_100) begin
        debug_4_12 = 1'b1;
      end else begin
        debug_4_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_100) begin
        debug_4_12 = 1'b1;
      end else begin
        debug_4_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_12 = 1'b0;
    if(when_ArraySlice_l165_101) begin
      if(when_ArraySlice_l166_101) begin
        debug_5_12 = 1'b1;
      end else begin
        debug_5_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_101) begin
        debug_5_12 = 1'b1;
      end else begin
        debug_5_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_12 = 1'b0;
    if(when_ArraySlice_l165_102) begin
      if(when_ArraySlice_l166_102) begin
        debug_6_12 = 1'b1;
      end else begin
        debug_6_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_102) begin
        debug_6_12 = 1'b1;
      end else begin
        debug_6_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_12 = 1'b0;
    if(when_ArraySlice_l165_103) begin
      if(when_ArraySlice_l166_103) begin
        debug_7_12 = 1'b1;
      end else begin
        debug_7_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_103) begin
        debug_7_12 = 1'b1;
      end else begin
        debug_7_12 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_96 = (_zz_when_ArraySlice_l165_96 <= selectWriteFifo);
  assign when_ArraySlice_l166_96 = (_zz_when_ArraySlice_l166_96 <= _zz_when_ArraySlice_l166_96_1);
  assign _zz_when_ArraySlice_l112_96 = (wReg % _zz__zz_when_ArraySlice_l112_96);
  assign when_ArraySlice_l112_96 = (_zz_when_ArraySlice_l112_96 != 6'h0);
  assign when_ArraySlice_l113_96 = (7'h40 <= _zz_when_ArraySlice_l113_96);
  always @(*) begin
    if(when_ArraySlice_l112_96) begin
      if(when_ArraySlice_l113_96) begin
        _zz_when_ArraySlice_l173_96 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_96 = (_zz__zz_when_ArraySlice_l173_96 - _zz__zz_when_ArraySlice_l173_96_3);
      end
    end else begin
      if(when_ArraySlice_l118_96) begin
        _zz_when_ArraySlice_l173_96 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_96 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_96 = (_zz_when_ArraySlice_l118_96 <= wReg);
  assign when_ArraySlice_l173_96 = (_zz_when_ArraySlice_l173_96_1 <= _zz_when_ArraySlice_l173_96_2);
  assign when_ArraySlice_l165_97 = (_zz_when_ArraySlice_l165_97 <= selectWriteFifo);
  assign when_ArraySlice_l166_97 = (_zz_when_ArraySlice_l166_97 <= _zz_when_ArraySlice_l166_97_1);
  assign _zz_when_ArraySlice_l112_97 = (wReg % _zz__zz_when_ArraySlice_l112_97);
  assign when_ArraySlice_l112_97 = (_zz_when_ArraySlice_l112_97 != 6'h0);
  assign when_ArraySlice_l113_97 = (7'h40 <= _zz_when_ArraySlice_l113_97);
  always @(*) begin
    if(when_ArraySlice_l112_97) begin
      if(when_ArraySlice_l113_97) begin
        _zz_when_ArraySlice_l173_97 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_97 = (_zz__zz_when_ArraySlice_l173_97 - _zz__zz_when_ArraySlice_l173_97_3);
      end
    end else begin
      if(when_ArraySlice_l118_97) begin
        _zz_when_ArraySlice_l173_97 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_97 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_97 = (_zz_when_ArraySlice_l118_97 <= wReg);
  assign when_ArraySlice_l173_97 = (_zz_when_ArraySlice_l173_97_1 <= _zz_when_ArraySlice_l173_97_3);
  assign when_ArraySlice_l165_98 = (_zz_when_ArraySlice_l165_98 <= selectWriteFifo);
  assign when_ArraySlice_l166_98 = (_zz_when_ArraySlice_l166_98 <= _zz_when_ArraySlice_l166_98_1);
  assign _zz_when_ArraySlice_l112_98 = (wReg % _zz__zz_when_ArraySlice_l112_98);
  assign when_ArraySlice_l112_98 = (_zz_when_ArraySlice_l112_98 != 6'h0);
  assign when_ArraySlice_l113_98 = (7'h40 <= _zz_when_ArraySlice_l113_98);
  always @(*) begin
    if(when_ArraySlice_l112_98) begin
      if(when_ArraySlice_l113_98) begin
        _zz_when_ArraySlice_l173_98 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_98 = (_zz__zz_when_ArraySlice_l173_98 - _zz__zz_when_ArraySlice_l173_98_3);
      end
    end else begin
      if(when_ArraySlice_l118_98) begin
        _zz_when_ArraySlice_l173_98 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_98 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_98 = (_zz_when_ArraySlice_l118_98 <= wReg);
  assign when_ArraySlice_l173_98 = (_zz_when_ArraySlice_l173_98_1 <= _zz_when_ArraySlice_l173_98_3);
  assign when_ArraySlice_l165_99 = (_zz_when_ArraySlice_l165_99 <= selectWriteFifo);
  assign when_ArraySlice_l166_99 = (_zz_when_ArraySlice_l166_99 <= _zz_when_ArraySlice_l166_99_1);
  assign _zz_when_ArraySlice_l112_99 = (wReg % _zz__zz_when_ArraySlice_l112_99);
  assign when_ArraySlice_l112_99 = (_zz_when_ArraySlice_l112_99 != 6'h0);
  assign when_ArraySlice_l113_99 = (7'h40 <= _zz_when_ArraySlice_l113_99);
  always @(*) begin
    if(when_ArraySlice_l112_99) begin
      if(when_ArraySlice_l113_99) begin
        _zz_when_ArraySlice_l173_99 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_99 = (_zz__zz_when_ArraySlice_l173_99 - _zz__zz_when_ArraySlice_l173_99_3);
      end
    end else begin
      if(when_ArraySlice_l118_99) begin
        _zz_when_ArraySlice_l173_99 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_99 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_99 = (_zz_when_ArraySlice_l118_99 <= wReg);
  assign when_ArraySlice_l173_99 = (_zz_when_ArraySlice_l173_99_1 <= _zz_when_ArraySlice_l173_99_3);
  assign when_ArraySlice_l165_100 = (_zz_when_ArraySlice_l165_100 <= selectWriteFifo);
  assign when_ArraySlice_l166_100 = (_zz_when_ArraySlice_l166_100 <= _zz_when_ArraySlice_l166_100_1);
  assign _zz_when_ArraySlice_l112_100 = (wReg % _zz__zz_when_ArraySlice_l112_100);
  assign when_ArraySlice_l112_100 = (_zz_when_ArraySlice_l112_100 != 6'h0);
  assign when_ArraySlice_l113_100 = (7'h40 <= _zz_when_ArraySlice_l113_100);
  always @(*) begin
    if(when_ArraySlice_l112_100) begin
      if(when_ArraySlice_l113_100) begin
        _zz_when_ArraySlice_l173_100 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_100 = (_zz__zz_when_ArraySlice_l173_100 - _zz__zz_when_ArraySlice_l173_100_3);
      end
    end else begin
      if(when_ArraySlice_l118_100) begin
        _zz_when_ArraySlice_l173_100 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_100 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_100 = (_zz_when_ArraySlice_l118_100 <= wReg);
  assign when_ArraySlice_l173_100 = (_zz_when_ArraySlice_l173_100_1 <= _zz_when_ArraySlice_l173_100_3);
  assign when_ArraySlice_l165_101 = (_zz_when_ArraySlice_l165_101 <= selectWriteFifo);
  assign when_ArraySlice_l166_101 = (_zz_when_ArraySlice_l166_101 <= _zz_when_ArraySlice_l166_101_2);
  assign _zz_when_ArraySlice_l112_101 = (wReg % _zz__zz_when_ArraySlice_l112_101);
  assign when_ArraySlice_l112_101 = (_zz_when_ArraySlice_l112_101 != 6'h0);
  assign when_ArraySlice_l113_101 = (7'h40 <= _zz_when_ArraySlice_l113_101);
  always @(*) begin
    if(when_ArraySlice_l112_101) begin
      if(when_ArraySlice_l113_101) begin
        _zz_when_ArraySlice_l173_101 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_101 = (_zz__zz_when_ArraySlice_l173_101 - _zz__zz_when_ArraySlice_l173_101_3);
      end
    end else begin
      if(when_ArraySlice_l118_101) begin
        _zz_when_ArraySlice_l173_101 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_101 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_101 = (_zz_when_ArraySlice_l118_101 <= wReg);
  assign when_ArraySlice_l173_101 = (_zz_when_ArraySlice_l173_101_1 <= _zz_when_ArraySlice_l173_101_3);
  assign when_ArraySlice_l165_102 = (_zz_when_ArraySlice_l165_102 <= selectWriteFifo);
  assign when_ArraySlice_l166_102 = (_zz_when_ArraySlice_l166_102 <= _zz_when_ArraySlice_l166_102_2);
  assign _zz_when_ArraySlice_l112_102 = (wReg % _zz__zz_when_ArraySlice_l112_102);
  assign when_ArraySlice_l112_102 = (_zz_when_ArraySlice_l112_102 != 6'h0);
  assign when_ArraySlice_l113_102 = (7'h40 <= _zz_when_ArraySlice_l113_102);
  always @(*) begin
    if(when_ArraySlice_l112_102) begin
      if(when_ArraySlice_l113_102) begin
        _zz_when_ArraySlice_l173_102 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_102 = (_zz__zz_when_ArraySlice_l173_102 - _zz__zz_when_ArraySlice_l173_102_3);
      end
    end else begin
      if(when_ArraySlice_l118_102) begin
        _zz_when_ArraySlice_l173_102 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_102 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_102 = (_zz_when_ArraySlice_l118_102 <= wReg);
  assign when_ArraySlice_l173_102 = (_zz_when_ArraySlice_l173_102_1 <= _zz_when_ArraySlice_l173_102_3);
  assign when_ArraySlice_l165_103 = (_zz_when_ArraySlice_l165_103 <= selectWriteFifo);
  assign when_ArraySlice_l166_103 = (_zz_when_ArraySlice_l166_103 <= _zz_when_ArraySlice_l166_103_2);
  assign _zz_when_ArraySlice_l112_103 = (wReg % _zz__zz_when_ArraySlice_l112_103);
  assign when_ArraySlice_l112_103 = (_zz_when_ArraySlice_l112_103 != 6'h0);
  assign when_ArraySlice_l113_103 = (7'h40 <= _zz_when_ArraySlice_l113_103);
  always @(*) begin
    if(when_ArraySlice_l112_103) begin
      if(when_ArraySlice_l113_103) begin
        _zz_when_ArraySlice_l173_103 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_103 = (_zz__zz_when_ArraySlice_l173_103 - _zz__zz_when_ArraySlice_l173_103_3);
      end
    end else begin
      if(when_ArraySlice_l118_103) begin
        _zz_when_ArraySlice_l173_103 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_103 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_103 = (_zz_when_ArraySlice_l118_103 <= wReg);
  assign when_ArraySlice_l173_103 = (_zz_when_ArraySlice_l173_103_1 <= _zz_when_ArraySlice_l173_103_3);
  assign when_ArraySlice_l444_3 = (! ((((((_zz_when_ArraySlice_l444_3_1 && _zz_when_ArraySlice_l444_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l444_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l444_3_4 && _zz_when_ArraySlice_l444_3_5) && (debug_4_12 == _zz_when_ArraySlice_l444_3_6)) && (debug_5_12 == 1'b1)) && (debug_6_12 == 1'b1)) && (debug_7_12 == 1'b1))));
  assign outputStreamArrayData_3_fire_5 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l448_3 = ((_zz_when_ArraySlice_l448_3_1 == 13'h0) && outputStreamArrayData_3_fire_5);
  assign when_ArraySlice_l434_3 = (allowPadding_3 && (wReg <= _zz_when_ArraySlice_l434_3));
  assign outputStreamArrayData_3_fire_6 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l455_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l455_3_1);
  assign when_ArraySlice_l373_4 = (_zz_when_ArraySlice_l373_4 < wReg);
  assign when_ArraySlice_l374_4 = ((! holdReadOp_4) && (_zz_when_ArraySlice_l374_4 != 7'h0));
  assign _zz_outputStreamArrayData_4_valid = (selectReadFifo_4 + _zz__zz_outputStreamArrayData_4_valid);
  assign _zz_7 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_4_valid);
  assign _zz_io_pop_ready_4 = outputStreamArrayData_4_ready;
  assign when_ArraySlice_l379_4 = (! holdReadOp_4);
  assign outputStreamArrayData_4_fire = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l380_4 = ((_zz_when_ArraySlice_l380_4_1 < _zz_when_ArraySlice_l380_4_3) && outputStreamArrayData_4_fire);
  assign when_ArraySlice_l381_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l381_4_1);
  assign when_ArraySlice_l384_4 = (_zz_when_ArraySlice_l384_4 == 13'h0);
  assign outputStreamArrayData_4_fire_1 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l389_4 = ((_zz_when_ArraySlice_l389_4_1 == _zz_when_ArraySlice_l389_4_4) && outputStreamArrayData_4_fire_1);
  assign when_ArraySlice_l390_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l390_4_1);
  assign _zz_when_ArraySlice_l94_12 = (hReg % _zz__zz_when_ArraySlice_l94_12);
  assign when_ArraySlice_l94_12 = (_zz_when_ArraySlice_l94_12 != 6'h0);
  assign when_ArraySlice_l95_12 = (7'h40 <= _zz_when_ArraySlice_l95_12);
  always @(*) begin
    if(when_ArraySlice_l94_12) begin
      if(when_ArraySlice_l95_12) begin
        _zz_when_ArraySlice_l392_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_4 = (_zz__zz_when_ArraySlice_l392_4 - _zz__zz_when_ArraySlice_l392_4_3);
      end
    end else begin
      if(when_ArraySlice_l99_12) begin
        _zz_when_ArraySlice_l392_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_4 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_12 = (_zz_when_ArraySlice_l99_12 <= hReg);
  assign when_ArraySlice_l392_4 = (_zz_when_ArraySlice_l392_4_1 < _zz_when_ArraySlice_l392_4_4);
  always @(*) begin
    debug_0_13 = 1'b0;
    if(when_ArraySlice_l165_104) begin
      if(when_ArraySlice_l166_104) begin
        debug_0_13 = 1'b1;
      end else begin
        debug_0_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_104) begin
        debug_0_13 = 1'b1;
      end else begin
        debug_0_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_13 = 1'b0;
    if(when_ArraySlice_l165_105) begin
      if(when_ArraySlice_l166_105) begin
        debug_1_13 = 1'b1;
      end else begin
        debug_1_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_105) begin
        debug_1_13 = 1'b1;
      end else begin
        debug_1_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_13 = 1'b0;
    if(when_ArraySlice_l165_106) begin
      if(when_ArraySlice_l166_106) begin
        debug_2_13 = 1'b1;
      end else begin
        debug_2_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_106) begin
        debug_2_13 = 1'b1;
      end else begin
        debug_2_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_13 = 1'b0;
    if(when_ArraySlice_l165_107) begin
      if(when_ArraySlice_l166_107) begin
        debug_3_13 = 1'b1;
      end else begin
        debug_3_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_107) begin
        debug_3_13 = 1'b1;
      end else begin
        debug_3_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_13 = 1'b0;
    if(when_ArraySlice_l165_108) begin
      if(when_ArraySlice_l166_108) begin
        debug_4_13 = 1'b1;
      end else begin
        debug_4_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_108) begin
        debug_4_13 = 1'b1;
      end else begin
        debug_4_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_13 = 1'b0;
    if(when_ArraySlice_l165_109) begin
      if(when_ArraySlice_l166_109) begin
        debug_5_13 = 1'b1;
      end else begin
        debug_5_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_109) begin
        debug_5_13 = 1'b1;
      end else begin
        debug_5_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_13 = 1'b0;
    if(when_ArraySlice_l165_110) begin
      if(when_ArraySlice_l166_110) begin
        debug_6_13 = 1'b1;
      end else begin
        debug_6_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_110) begin
        debug_6_13 = 1'b1;
      end else begin
        debug_6_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_13 = 1'b0;
    if(when_ArraySlice_l165_111) begin
      if(when_ArraySlice_l166_111) begin
        debug_7_13 = 1'b1;
      end else begin
        debug_7_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_111) begin
        debug_7_13 = 1'b1;
      end else begin
        debug_7_13 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_104 = (_zz_when_ArraySlice_l165_104 <= selectWriteFifo);
  assign when_ArraySlice_l166_104 = (_zz_when_ArraySlice_l166_104 <= _zz_when_ArraySlice_l166_104_1);
  assign _zz_when_ArraySlice_l112_104 = (wReg % _zz__zz_when_ArraySlice_l112_104);
  assign when_ArraySlice_l112_104 = (_zz_when_ArraySlice_l112_104 != 6'h0);
  assign when_ArraySlice_l113_104 = (7'h40 <= _zz_when_ArraySlice_l113_104);
  always @(*) begin
    if(when_ArraySlice_l112_104) begin
      if(when_ArraySlice_l113_104) begin
        _zz_when_ArraySlice_l173_104 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_104 = (_zz__zz_when_ArraySlice_l173_104 - _zz__zz_when_ArraySlice_l173_104_3);
      end
    end else begin
      if(when_ArraySlice_l118_104) begin
        _zz_when_ArraySlice_l173_104 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_104 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_104 = (_zz_when_ArraySlice_l118_104 <= wReg);
  assign when_ArraySlice_l173_104 = (_zz_when_ArraySlice_l173_104_1 <= _zz_when_ArraySlice_l173_104_2);
  assign when_ArraySlice_l165_105 = (_zz_when_ArraySlice_l165_105 <= selectWriteFifo);
  assign when_ArraySlice_l166_105 = (_zz_when_ArraySlice_l166_105 <= _zz_when_ArraySlice_l166_105_1);
  assign _zz_when_ArraySlice_l112_105 = (wReg % _zz__zz_when_ArraySlice_l112_105);
  assign when_ArraySlice_l112_105 = (_zz_when_ArraySlice_l112_105 != 6'h0);
  assign when_ArraySlice_l113_105 = (7'h40 <= _zz_when_ArraySlice_l113_105);
  always @(*) begin
    if(when_ArraySlice_l112_105) begin
      if(when_ArraySlice_l113_105) begin
        _zz_when_ArraySlice_l173_105 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_105 = (_zz__zz_when_ArraySlice_l173_105 - _zz__zz_when_ArraySlice_l173_105_3);
      end
    end else begin
      if(when_ArraySlice_l118_105) begin
        _zz_when_ArraySlice_l173_105 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_105 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_105 = (_zz_when_ArraySlice_l118_105 <= wReg);
  assign when_ArraySlice_l173_105 = (_zz_when_ArraySlice_l173_105_1 <= _zz_when_ArraySlice_l173_105_3);
  assign when_ArraySlice_l165_106 = (_zz_when_ArraySlice_l165_106 <= selectWriteFifo);
  assign when_ArraySlice_l166_106 = (_zz_when_ArraySlice_l166_106 <= _zz_when_ArraySlice_l166_106_1);
  assign _zz_when_ArraySlice_l112_106 = (wReg % _zz__zz_when_ArraySlice_l112_106);
  assign when_ArraySlice_l112_106 = (_zz_when_ArraySlice_l112_106 != 6'h0);
  assign when_ArraySlice_l113_106 = (7'h40 <= _zz_when_ArraySlice_l113_106);
  always @(*) begin
    if(when_ArraySlice_l112_106) begin
      if(when_ArraySlice_l113_106) begin
        _zz_when_ArraySlice_l173_106 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_106 = (_zz__zz_when_ArraySlice_l173_106 - _zz__zz_when_ArraySlice_l173_106_3);
      end
    end else begin
      if(when_ArraySlice_l118_106) begin
        _zz_when_ArraySlice_l173_106 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_106 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_106 = (_zz_when_ArraySlice_l118_106 <= wReg);
  assign when_ArraySlice_l173_106 = (_zz_when_ArraySlice_l173_106_1 <= _zz_when_ArraySlice_l173_106_3);
  assign when_ArraySlice_l165_107 = (_zz_when_ArraySlice_l165_107 <= selectWriteFifo);
  assign when_ArraySlice_l166_107 = (_zz_when_ArraySlice_l166_107 <= _zz_when_ArraySlice_l166_107_1);
  assign _zz_when_ArraySlice_l112_107 = (wReg % _zz__zz_when_ArraySlice_l112_107);
  assign when_ArraySlice_l112_107 = (_zz_when_ArraySlice_l112_107 != 6'h0);
  assign when_ArraySlice_l113_107 = (7'h40 <= _zz_when_ArraySlice_l113_107);
  always @(*) begin
    if(when_ArraySlice_l112_107) begin
      if(when_ArraySlice_l113_107) begin
        _zz_when_ArraySlice_l173_107 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_107 = (_zz__zz_when_ArraySlice_l173_107 - _zz__zz_when_ArraySlice_l173_107_3);
      end
    end else begin
      if(when_ArraySlice_l118_107) begin
        _zz_when_ArraySlice_l173_107 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_107 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_107 = (_zz_when_ArraySlice_l118_107 <= wReg);
  assign when_ArraySlice_l173_107 = (_zz_when_ArraySlice_l173_107_1 <= _zz_when_ArraySlice_l173_107_3);
  assign when_ArraySlice_l165_108 = (_zz_when_ArraySlice_l165_108 <= selectWriteFifo);
  assign when_ArraySlice_l166_108 = (_zz_when_ArraySlice_l166_108 <= _zz_when_ArraySlice_l166_108_1);
  assign _zz_when_ArraySlice_l112_108 = (wReg % _zz__zz_when_ArraySlice_l112_108);
  assign when_ArraySlice_l112_108 = (_zz_when_ArraySlice_l112_108 != 6'h0);
  assign when_ArraySlice_l113_108 = (7'h40 <= _zz_when_ArraySlice_l113_108);
  always @(*) begin
    if(when_ArraySlice_l112_108) begin
      if(when_ArraySlice_l113_108) begin
        _zz_when_ArraySlice_l173_108 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_108 = (_zz__zz_when_ArraySlice_l173_108 - _zz__zz_when_ArraySlice_l173_108_3);
      end
    end else begin
      if(when_ArraySlice_l118_108) begin
        _zz_when_ArraySlice_l173_108 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_108 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_108 = (_zz_when_ArraySlice_l118_108 <= wReg);
  assign when_ArraySlice_l173_108 = (_zz_when_ArraySlice_l173_108_1 <= _zz_when_ArraySlice_l173_108_3);
  assign when_ArraySlice_l165_109 = (_zz_when_ArraySlice_l165_109 <= selectWriteFifo);
  assign when_ArraySlice_l166_109 = (_zz_when_ArraySlice_l166_109 <= _zz_when_ArraySlice_l166_109_2);
  assign _zz_when_ArraySlice_l112_109 = (wReg % _zz__zz_when_ArraySlice_l112_109);
  assign when_ArraySlice_l112_109 = (_zz_when_ArraySlice_l112_109 != 6'h0);
  assign when_ArraySlice_l113_109 = (7'h40 <= _zz_when_ArraySlice_l113_109);
  always @(*) begin
    if(when_ArraySlice_l112_109) begin
      if(when_ArraySlice_l113_109) begin
        _zz_when_ArraySlice_l173_109 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_109 = (_zz__zz_when_ArraySlice_l173_109 - _zz__zz_when_ArraySlice_l173_109_3);
      end
    end else begin
      if(when_ArraySlice_l118_109) begin
        _zz_when_ArraySlice_l173_109 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_109 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_109 = (_zz_when_ArraySlice_l118_109 <= wReg);
  assign when_ArraySlice_l173_109 = (_zz_when_ArraySlice_l173_109_1 <= _zz_when_ArraySlice_l173_109_3);
  assign when_ArraySlice_l165_110 = (_zz_when_ArraySlice_l165_110 <= selectWriteFifo);
  assign when_ArraySlice_l166_110 = (_zz_when_ArraySlice_l166_110 <= _zz_when_ArraySlice_l166_110_2);
  assign _zz_when_ArraySlice_l112_110 = (wReg % _zz__zz_when_ArraySlice_l112_110);
  assign when_ArraySlice_l112_110 = (_zz_when_ArraySlice_l112_110 != 6'h0);
  assign when_ArraySlice_l113_110 = (7'h40 <= _zz_when_ArraySlice_l113_110);
  always @(*) begin
    if(when_ArraySlice_l112_110) begin
      if(when_ArraySlice_l113_110) begin
        _zz_when_ArraySlice_l173_110 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_110 = (_zz__zz_when_ArraySlice_l173_110 - _zz__zz_when_ArraySlice_l173_110_3);
      end
    end else begin
      if(when_ArraySlice_l118_110) begin
        _zz_when_ArraySlice_l173_110 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_110 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_110 = (_zz_when_ArraySlice_l118_110 <= wReg);
  assign when_ArraySlice_l173_110 = (_zz_when_ArraySlice_l173_110_1 <= _zz_when_ArraySlice_l173_110_3);
  assign when_ArraySlice_l165_111 = (_zz_when_ArraySlice_l165_111 <= selectWriteFifo);
  assign when_ArraySlice_l166_111 = (_zz_when_ArraySlice_l166_111 <= _zz_when_ArraySlice_l166_111_2);
  assign _zz_when_ArraySlice_l112_111 = (wReg % _zz__zz_when_ArraySlice_l112_111);
  assign when_ArraySlice_l112_111 = (_zz_when_ArraySlice_l112_111 != 6'h0);
  assign when_ArraySlice_l113_111 = (7'h40 <= _zz_when_ArraySlice_l113_111);
  always @(*) begin
    if(when_ArraySlice_l112_111) begin
      if(when_ArraySlice_l113_111) begin
        _zz_when_ArraySlice_l173_111 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_111 = (_zz__zz_when_ArraySlice_l173_111 - _zz__zz_when_ArraySlice_l173_111_3);
      end
    end else begin
      if(when_ArraySlice_l118_111) begin
        _zz_when_ArraySlice_l173_111 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_111 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_111 = (_zz_when_ArraySlice_l118_111 <= wReg);
  assign when_ArraySlice_l173_111 = (_zz_when_ArraySlice_l173_111_1 <= _zz_when_ArraySlice_l173_111_3);
  assign when_ArraySlice_l398_4 = (! ((((((_zz_when_ArraySlice_l398_4_1 && _zz_when_ArraySlice_l398_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l398_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l398_4_4 && _zz_when_ArraySlice_l398_4_5) && (debug_4_13 == _zz_when_ArraySlice_l398_4_6)) && (debug_5_13 == 1'b1)) && (debug_6_13 == 1'b1)) && (debug_7_13 == 1'b1))));
  assign when_ArraySlice_l401_4 = (wReg <= _zz_when_ArraySlice_l401_4_1);
  assign when_ArraySlice_l405_4 = (_zz_when_ArraySlice_l405_4 == 13'h0);
  assign when_ArraySlice_l409_4 = (_zz_when_ArraySlice_l409_4 == 7'h0);
  assign outputStreamArrayData_4_fire_2 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l410_4 = ((handshakeTimes_4_value == _zz_when_ArraySlice_l410_4_1) && outputStreamArrayData_4_fire_2);
  assign _zz_when_ArraySlice_l94_13 = (hReg % _zz__zz_when_ArraySlice_l94_13);
  assign when_ArraySlice_l94_13 = (_zz_when_ArraySlice_l94_13 != 6'h0);
  assign when_ArraySlice_l95_13 = (7'h40 <= _zz_when_ArraySlice_l95_13);
  always @(*) begin
    if(when_ArraySlice_l94_13) begin
      if(when_ArraySlice_l95_13) begin
        _zz_when_ArraySlice_l412_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_4 = (_zz__zz_when_ArraySlice_l412_4 - _zz__zz_when_ArraySlice_l412_4_3);
      end
    end else begin
      if(when_ArraySlice_l99_13) begin
        _zz_when_ArraySlice_l412_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_4 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_13 = (_zz_when_ArraySlice_l99_13 <= hReg);
  assign when_ArraySlice_l412_4 = (_zz_when_ArraySlice_l412_4_1 < _zz_when_ArraySlice_l412_4_4);
  always @(*) begin
    debug_0_14 = 1'b0;
    if(when_ArraySlice_l165_112) begin
      if(when_ArraySlice_l166_112) begin
        debug_0_14 = 1'b1;
      end else begin
        debug_0_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_112) begin
        debug_0_14 = 1'b1;
      end else begin
        debug_0_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_14 = 1'b0;
    if(when_ArraySlice_l165_113) begin
      if(when_ArraySlice_l166_113) begin
        debug_1_14 = 1'b1;
      end else begin
        debug_1_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_113) begin
        debug_1_14 = 1'b1;
      end else begin
        debug_1_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_14 = 1'b0;
    if(when_ArraySlice_l165_114) begin
      if(when_ArraySlice_l166_114) begin
        debug_2_14 = 1'b1;
      end else begin
        debug_2_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_114) begin
        debug_2_14 = 1'b1;
      end else begin
        debug_2_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_14 = 1'b0;
    if(when_ArraySlice_l165_115) begin
      if(when_ArraySlice_l166_115) begin
        debug_3_14 = 1'b1;
      end else begin
        debug_3_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_115) begin
        debug_3_14 = 1'b1;
      end else begin
        debug_3_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_14 = 1'b0;
    if(when_ArraySlice_l165_116) begin
      if(when_ArraySlice_l166_116) begin
        debug_4_14 = 1'b1;
      end else begin
        debug_4_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_116) begin
        debug_4_14 = 1'b1;
      end else begin
        debug_4_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_14 = 1'b0;
    if(when_ArraySlice_l165_117) begin
      if(when_ArraySlice_l166_117) begin
        debug_5_14 = 1'b1;
      end else begin
        debug_5_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_117) begin
        debug_5_14 = 1'b1;
      end else begin
        debug_5_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_14 = 1'b0;
    if(when_ArraySlice_l165_118) begin
      if(when_ArraySlice_l166_118) begin
        debug_6_14 = 1'b1;
      end else begin
        debug_6_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_118) begin
        debug_6_14 = 1'b1;
      end else begin
        debug_6_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_14 = 1'b0;
    if(when_ArraySlice_l165_119) begin
      if(when_ArraySlice_l166_119) begin
        debug_7_14 = 1'b1;
      end else begin
        debug_7_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_119) begin
        debug_7_14 = 1'b1;
      end else begin
        debug_7_14 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_112 = (_zz_when_ArraySlice_l165_112 <= selectWriteFifo);
  assign when_ArraySlice_l166_112 = (_zz_when_ArraySlice_l166_112 <= _zz_when_ArraySlice_l166_112_1);
  assign _zz_when_ArraySlice_l112_112 = (wReg % _zz__zz_when_ArraySlice_l112_112);
  assign when_ArraySlice_l112_112 = (_zz_when_ArraySlice_l112_112 != 6'h0);
  assign when_ArraySlice_l113_112 = (7'h40 <= _zz_when_ArraySlice_l113_112);
  always @(*) begin
    if(when_ArraySlice_l112_112) begin
      if(when_ArraySlice_l113_112) begin
        _zz_when_ArraySlice_l173_112 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_112 = (_zz__zz_when_ArraySlice_l173_112 - _zz__zz_when_ArraySlice_l173_112_3);
      end
    end else begin
      if(when_ArraySlice_l118_112) begin
        _zz_when_ArraySlice_l173_112 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_112 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_112 = (_zz_when_ArraySlice_l118_112 <= wReg);
  assign when_ArraySlice_l173_112 = (_zz_when_ArraySlice_l173_112_1 <= _zz_when_ArraySlice_l173_112_2);
  assign when_ArraySlice_l165_113 = (_zz_when_ArraySlice_l165_113 <= selectWriteFifo);
  assign when_ArraySlice_l166_113 = (_zz_when_ArraySlice_l166_113 <= _zz_when_ArraySlice_l166_113_1);
  assign _zz_when_ArraySlice_l112_113 = (wReg % _zz__zz_when_ArraySlice_l112_113);
  assign when_ArraySlice_l112_113 = (_zz_when_ArraySlice_l112_113 != 6'h0);
  assign when_ArraySlice_l113_113 = (7'h40 <= _zz_when_ArraySlice_l113_113);
  always @(*) begin
    if(when_ArraySlice_l112_113) begin
      if(when_ArraySlice_l113_113) begin
        _zz_when_ArraySlice_l173_113 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_113 = (_zz__zz_when_ArraySlice_l173_113 - _zz__zz_when_ArraySlice_l173_113_3);
      end
    end else begin
      if(when_ArraySlice_l118_113) begin
        _zz_when_ArraySlice_l173_113 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_113 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_113 = (_zz_when_ArraySlice_l118_113 <= wReg);
  assign when_ArraySlice_l173_113 = (_zz_when_ArraySlice_l173_113_1 <= _zz_when_ArraySlice_l173_113_3);
  assign when_ArraySlice_l165_114 = (_zz_when_ArraySlice_l165_114 <= selectWriteFifo);
  assign when_ArraySlice_l166_114 = (_zz_when_ArraySlice_l166_114 <= _zz_when_ArraySlice_l166_114_1);
  assign _zz_when_ArraySlice_l112_114 = (wReg % _zz__zz_when_ArraySlice_l112_114);
  assign when_ArraySlice_l112_114 = (_zz_when_ArraySlice_l112_114 != 6'h0);
  assign when_ArraySlice_l113_114 = (7'h40 <= _zz_when_ArraySlice_l113_114);
  always @(*) begin
    if(when_ArraySlice_l112_114) begin
      if(when_ArraySlice_l113_114) begin
        _zz_when_ArraySlice_l173_114 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_114 = (_zz__zz_when_ArraySlice_l173_114 - _zz__zz_when_ArraySlice_l173_114_3);
      end
    end else begin
      if(when_ArraySlice_l118_114) begin
        _zz_when_ArraySlice_l173_114 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_114 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_114 = (_zz_when_ArraySlice_l118_114 <= wReg);
  assign when_ArraySlice_l173_114 = (_zz_when_ArraySlice_l173_114_1 <= _zz_when_ArraySlice_l173_114_3);
  assign when_ArraySlice_l165_115 = (_zz_when_ArraySlice_l165_115 <= selectWriteFifo);
  assign when_ArraySlice_l166_115 = (_zz_when_ArraySlice_l166_115 <= _zz_when_ArraySlice_l166_115_1);
  assign _zz_when_ArraySlice_l112_115 = (wReg % _zz__zz_when_ArraySlice_l112_115);
  assign when_ArraySlice_l112_115 = (_zz_when_ArraySlice_l112_115 != 6'h0);
  assign when_ArraySlice_l113_115 = (7'h40 <= _zz_when_ArraySlice_l113_115);
  always @(*) begin
    if(when_ArraySlice_l112_115) begin
      if(when_ArraySlice_l113_115) begin
        _zz_when_ArraySlice_l173_115 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_115 = (_zz__zz_when_ArraySlice_l173_115 - _zz__zz_when_ArraySlice_l173_115_3);
      end
    end else begin
      if(when_ArraySlice_l118_115) begin
        _zz_when_ArraySlice_l173_115 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_115 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_115 = (_zz_when_ArraySlice_l118_115 <= wReg);
  assign when_ArraySlice_l173_115 = (_zz_when_ArraySlice_l173_115_1 <= _zz_when_ArraySlice_l173_115_3);
  assign when_ArraySlice_l165_116 = (_zz_when_ArraySlice_l165_116 <= selectWriteFifo);
  assign when_ArraySlice_l166_116 = (_zz_when_ArraySlice_l166_116 <= _zz_when_ArraySlice_l166_116_1);
  assign _zz_when_ArraySlice_l112_116 = (wReg % _zz__zz_when_ArraySlice_l112_116);
  assign when_ArraySlice_l112_116 = (_zz_when_ArraySlice_l112_116 != 6'h0);
  assign when_ArraySlice_l113_116 = (7'h40 <= _zz_when_ArraySlice_l113_116);
  always @(*) begin
    if(when_ArraySlice_l112_116) begin
      if(when_ArraySlice_l113_116) begin
        _zz_when_ArraySlice_l173_116 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_116 = (_zz__zz_when_ArraySlice_l173_116 - _zz__zz_when_ArraySlice_l173_116_3);
      end
    end else begin
      if(when_ArraySlice_l118_116) begin
        _zz_when_ArraySlice_l173_116 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_116 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_116 = (_zz_when_ArraySlice_l118_116 <= wReg);
  assign when_ArraySlice_l173_116 = (_zz_when_ArraySlice_l173_116_1 <= _zz_when_ArraySlice_l173_116_3);
  assign when_ArraySlice_l165_117 = (_zz_when_ArraySlice_l165_117 <= selectWriteFifo);
  assign when_ArraySlice_l166_117 = (_zz_when_ArraySlice_l166_117 <= _zz_when_ArraySlice_l166_117_2);
  assign _zz_when_ArraySlice_l112_117 = (wReg % _zz__zz_when_ArraySlice_l112_117);
  assign when_ArraySlice_l112_117 = (_zz_when_ArraySlice_l112_117 != 6'h0);
  assign when_ArraySlice_l113_117 = (7'h40 <= _zz_when_ArraySlice_l113_117);
  always @(*) begin
    if(when_ArraySlice_l112_117) begin
      if(when_ArraySlice_l113_117) begin
        _zz_when_ArraySlice_l173_117 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_117 = (_zz__zz_when_ArraySlice_l173_117 - _zz__zz_when_ArraySlice_l173_117_3);
      end
    end else begin
      if(when_ArraySlice_l118_117) begin
        _zz_when_ArraySlice_l173_117 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_117 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_117 = (_zz_when_ArraySlice_l118_117 <= wReg);
  assign when_ArraySlice_l173_117 = (_zz_when_ArraySlice_l173_117_1 <= _zz_when_ArraySlice_l173_117_3);
  assign when_ArraySlice_l165_118 = (_zz_when_ArraySlice_l165_118 <= selectWriteFifo);
  assign when_ArraySlice_l166_118 = (_zz_when_ArraySlice_l166_118 <= _zz_when_ArraySlice_l166_118_2);
  assign _zz_when_ArraySlice_l112_118 = (wReg % _zz__zz_when_ArraySlice_l112_118);
  assign when_ArraySlice_l112_118 = (_zz_when_ArraySlice_l112_118 != 6'h0);
  assign when_ArraySlice_l113_118 = (7'h40 <= _zz_when_ArraySlice_l113_118);
  always @(*) begin
    if(when_ArraySlice_l112_118) begin
      if(when_ArraySlice_l113_118) begin
        _zz_when_ArraySlice_l173_118 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_118 = (_zz__zz_when_ArraySlice_l173_118 - _zz__zz_when_ArraySlice_l173_118_3);
      end
    end else begin
      if(when_ArraySlice_l118_118) begin
        _zz_when_ArraySlice_l173_118 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_118 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_118 = (_zz_when_ArraySlice_l118_118 <= wReg);
  assign when_ArraySlice_l173_118 = (_zz_when_ArraySlice_l173_118_1 <= _zz_when_ArraySlice_l173_118_3);
  assign when_ArraySlice_l165_119 = (_zz_when_ArraySlice_l165_119 <= selectWriteFifo);
  assign when_ArraySlice_l166_119 = (_zz_when_ArraySlice_l166_119 <= _zz_when_ArraySlice_l166_119_2);
  assign _zz_when_ArraySlice_l112_119 = (wReg % _zz__zz_when_ArraySlice_l112_119);
  assign when_ArraySlice_l112_119 = (_zz_when_ArraySlice_l112_119 != 6'h0);
  assign when_ArraySlice_l113_119 = (7'h40 <= _zz_when_ArraySlice_l113_119);
  always @(*) begin
    if(when_ArraySlice_l112_119) begin
      if(when_ArraySlice_l113_119) begin
        _zz_when_ArraySlice_l173_119 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_119 = (_zz__zz_when_ArraySlice_l173_119 - _zz__zz_when_ArraySlice_l173_119_3);
      end
    end else begin
      if(when_ArraySlice_l118_119) begin
        _zz_when_ArraySlice_l173_119 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_119 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_119 = (_zz_when_ArraySlice_l118_119 <= wReg);
  assign when_ArraySlice_l173_119 = (_zz_when_ArraySlice_l173_119_1 <= _zz_when_ArraySlice_l173_119_3);
  assign when_ArraySlice_l418_4 = (! ((((((_zz_when_ArraySlice_l418_4_1 && _zz_when_ArraySlice_l418_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l418_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l418_4_4 && _zz_when_ArraySlice_l418_4_5) && (debug_4_14 == _zz_when_ArraySlice_l418_4_6)) && (debug_5_14 == 1'b1)) && (debug_6_14 == 1'b1)) && (debug_7_14 == 1'b1))));
  assign when_ArraySlice_l421_4 = (wReg <= _zz_when_ArraySlice_l421_4_1);
  assign outputStreamArrayData_4_fire_3 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l425_4 = ((_zz_when_ArraySlice_l425_4 == 13'h0) && outputStreamArrayData_4_fire_3);
  assign outputStreamArrayData_4_fire_4 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l436_4 = ((handshakeTimes_4_value == _zz_when_ArraySlice_l436_4_1) && outputStreamArrayData_4_fire_4);
  assign _zz_when_ArraySlice_l94_14 = (hReg % _zz__zz_when_ArraySlice_l94_14);
  assign when_ArraySlice_l94_14 = (_zz_when_ArraySlice_l94_14 != 6'h0);
  assign when_ArraySlice_l95_14 = (7'h40 <= _zz_when_ArraySlice_l95_14);
  always @(*) begin
    if(when_ArraySlice_l94_14) begin
      if(when_ArraySlice_l95_14) begin
        _zz_when_ArraySlice_l437_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_4 = (_zz__zz_when_ArraySlice_l437_4 - _zz__zz_when_ArraySlice_l437_4_3);
      end
    end else begin
      if(when_ArraySlice_l99_14) begin
        _zz_when_ArraySlice_l437_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_4 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_14 = (_zz_when_ArraySlice_l99_14 <= hReg);
  assign when_ArraySlice_l437_4 = (_zz_when_ArraySlice_l437_4_1 < _zz_when_ArraySlice_l437_4_4);
  always @(*) begin
    debug_0_15 = 1'b0;
    if(when_ArraySlice_l165_120) begin
      if(when_ArraySlice_l166_120) begin
        debug_0_15 = 1'b1;
      end else begin
        debug_0_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_120) begin
        debug_0_15 = 1'b1;
      end else begin
        debug_0_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_15 = 1'b0;
    if(when_ArraySlice_l165_121) begin
      if(when_ArraySlice_l166_121) begin
        debug_1_15 = 1'b1;
      end else begin
        debug_1_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_121) begin
        debug_1_15 = 1'b1;
      end else begin
        debug_1_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_15 = 1'b0;
    if(when_ArraySlice_l165_122) begin
      if(when_ArraySlice_l166_122) begin
        debug_2_15 = 1'b1;
      end else begin
        debug_2_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_122) begin
        debug_2_15 = 1'b1;
      end else begin
        debug_2_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_15 = 1'b0;
    if(when_ArraySlice_l165_123) begin
      if(when_ArraySlice_l166_123) begin
        debug_3_15 = 1'b1;
      end else begin
        debug_3_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_123) begin
        debug_3_15 = 1'b1;
      end else begin
        debug_3_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_15 = 1'b0;
    if(when_ArraySlice_l165_124) begin
      if(when_ArraySlice_l166_124) begin
        debug_4_15 = 1'b1;
      end else begin
        debug_4_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_124) begin
        debug_4_15 = 1'b1;
      end else begin
        debug_4_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_15 = 1'b0;
    if(when_ArraySlice_l165_125) begin
      if(when_ArraySlice_l166_125) begin
        debug_5_15 = 1'b1;
      end else begin
        debug_5_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_125) begin
        debug_5_15 = 1'b1;
      end else begin
        debug_5_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_15 = 1'b0;
    if(when_ArraySlice_l165_126) begin
      if(when_ArraySlice_l166_126) begin
        debug_6_15 = 1'b1;
      end else begin
        debug_6_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_126) begin
        debug_6_15 = 1'b1;
      end else begin
        debug_6_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_15 = 1'b0;
    if(when_ArraySlice_l165_127) begin
      if(when_ArraySlice_l166_127) begin
        debug_7_15 = 1'b1;
      end else begin
        debug_7_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_127) begin
        debug_7_15 = 1'b1;
      end else begin
        debug_7_15 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_120 = (_zz_when_ArraySlice_l165_120 <= selectWriteFifo);
  assign when_ArraySlice_l166_120 = (_zz_when_ArraySlice_l166_120 <= _zz_when_ArraySlice_l166_120_1);
  assign _zz_when_ArraySlice_l112_120 = (wReg % _zz__zz_when_ArraySlice_l112_120);
  assign when_ArraySlice_l112_120 = (_zz_when_ArraySlice_l112_120 != 6'h0);
  assign when_ArraySlice_l113_120 = (7'h40 <= _zz_when_ArraySlice_l113_120);
  always @(*) begin
    if(when_ArraySlice_l112_120) begin
      if(when_ArraySlice_l113_120) begin
        _zz_when_ArraySlice_l173_120 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_120 = (_zz__zz_when_ArraySlice_l173_120 - _zz__zz_when_ArraySlice_l173_120_3);
      end
    end else begin
      if(when_ArraySlice_l118_120) begin
        _zz_when_ArraySlice_l173_120 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_120 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_120 = (_zz_when_ArraySlice_l118_120 <= wReg);
  assign when_ArraySlice_l173_120 = (_zz_when_ArraySlice_l173_120_1 <= _zz_when_ArraySlice_l173_120_2);
  assign when_ArraySlice_l165_121 = (_zz_when_ArraySlice_l165_121 <= selectWriteFifo);
  assign when_ArraySlice_l166_121 = (_zz_when_ArraySlice_l166_121 <= _zz_when_ArraySlice_l166_121_1);
  assign _zz_when_ArraySlice_l112_121 = (wReg % _zz__zz_when_ArraySlice_l112_121);
  assign when_ArraySlice_l112_121 = (_zz_when_ArraySlice_l112_121 != 6'h0);
  assign when_ArraySlice_l113_121 = (7'h40 <= _zz_when_ArraySlice_l113_121);
  always @(*) begin
    if(when_ArraySlice_l112_121) begin
      if(when_ArraySlice_l113_121) begin
        _zz_when_ArraySlice_l173_121 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_121 = (_zz__zz_when_ArraySlice_l173_121 - _zz__zz_when_ArraySlice_l173_121_3);
      end
    end else begin
      if(when_ArraySlice_l118_121) begin
        _zz_when_ArraySlice_l173_121 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_121 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_121 = (_zz_when_ArraySlice_l118_121 <= wReg);
  assign when_ArraySlice_l173_121 = (_zz_when_ArraySlice_l173_121_1 <= _zz_when_ArraySlice_l173_121_3);
  assign when_ArraySlice_l165_122 = (_zz_when_ArraySlice_l165_122 <= selectWriteFifo);
  assign when_ArraySlice_l166_122 = (_zz_when_ArraySlice_l166_122 <= _zz_when_ArraySlice_l166_122_1);
  assign _zz_when_ArraySlice_l112_122 = (wReg % _zz__zz_when_ArraySlice_l112_122);
  assign when_ArraySlice_l112_122 = (_zz_when_ArraySlice_l112_122 != 6'h0);
  assign when_ArraySlice_l113_122 = (7'h40 <= _zz_when_ArraySlice_l113_122);
  always @(*) begin
    if(when_ArraySlice_l112_122) begin
      if(when_ArraySlice_l113_122) begin
        _zz_when_ArraySlice_l173_122 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_122 = (_zz__zz_when_ArraySlice_l173_122 - _zz__zz_when_ArraySlice_l173_122_3);
      end
    end else begin
      if(when_ArraySlice_l118_122) begin
        _zz_when_ArraySlice_l173_122 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_122 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_122 = (_zz_when_ArraySlice_l118_122 <= wReg);
  assign when_ArraySlice_l173_122 = (_zz_when_ArraySlice_l173_122_1 <= _zz_when_ArraySlice_l173_122_3);
  assign when_ArraySlice_l165_123 = (_zz_when_ArraySlice_l165_123 <= selectWriteFifo);
  assign when_ArraySlice_l166_123 = (_zz_when_ArraySlice_l166_123 <= _zz_when_ArraySlice_l166_123_1);
  assign _zz_when_ArraySlice_l112_123 = (wReg % _zz__zz_when_ArraySlice_l112_123);
  assign when_ArraySlice_l112_123 = (_zz_when_ArraySlice_l112_123 != 6'h0);
  assign when_ArraySlice_l113_123 = (7'h40 <= _zz_when_ArraySlice_l113_123);
  always @(*) begin
    if(when_ArraySlice_l112_123) begin
      if(when_ArraySlice_l113_123) begin
        _zz_when_ArraySlice_l173_123 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_123 = (_zz__zz_when_ArraySlice_l173_123 - _zz__zz_when_ArraySlice_l173_123_3);
      end
    end else begin
      if(when_ArraySlice_l118_123) begin
        _zz_when_ArraySlice_l173_123 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_123 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_123 = (_zz_when_ArraySlice_l118_123 <= wReg);
  assign when_ArraySlice_l173_123 = (_zz_when_ArraySlice_l173_123_1 <= _zz_when_ArraySlice_l173_123_3);
  assign when_ArraySlice_l165_124 = (_zz_when_ArraySlice_l165_124 <= selectWriteFifo);
  assign when_ArraySlice_l166_124 = (_zz_when_ArraySlice_l166_124 <= _zz_when_ArraySlice_l166_124_1);
  assign _zz_when_ArraySlice_l112_124 = (wReg % _zz__zz_when_ArraySlice_l112_124);
  assign when_ArraySlice_l112_124 = (_zz_when_ArraySlice_l112_124 != 6'h0);
  assign when_ArraySlice_l113_124 = (7'h40 <= _zz_when_ArraySlice_l113_124);
  always @(*) begin
    if(when_ArraySlice_l112_124) begin
      if(when_ArraySlice_l113_124) begin
        _zz_when_ArraySlice_l173_124 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_124 = (_zz__zz_when_ArraySlice_l173_124 - _zz__zz_when_ArraySlice_l173_124_3);
      end
    end else begin
      if(when_ArraySlice_l118_124) begin
        _zz_when_ArraySlice_l173_124 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_124 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_124 = (_zz_when_ArraySlice_l118_124 <= wReg);
  assign when_ArraySlice_l173_124 = (_zz_when_ArraySlice_l173_124_1 <= _zz_when_ArraySlice_l173_124_3);
  assign when_ArraySlice_l165_125 = (_zz_when_ArraySlice_l165_125 <= selectWriteFifo);
  assign when_ArraySlice_l166_125 = (_zz_when_ArraySlice_l166_125 <= _zz_when_ArraySlice_l166_125_2);
  assign _zz_when_ArraySlice_l112_125 = (wReg % _zz__zz_when_ArraySlice_l112_125);
  assign when_ArraySlice_l112_125 = (_zz_when_ArraySlice_l112_125 != 6'h0);
  assign when_ArraySlice_l113_125 = (7'h40 <= _zz_when_ArraySlice_l113_125);
  always @(*) begin
    if(when_ArraySlice_l112_125) begin
      if(when_ArraySlice_l113_125) begin
        _zz_when_ArraySlice_l173_125 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_125 = (_zz__zz_when_ArraySlice_l173_125 - _zz__zz_when_ArraySlice_l173_125_3);
      end
    end else begin
      if(when_ArraySlice_l118_125) begin
        _zz_when_ArraySlice_l173_125 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_125 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_125 = (_zz_when_ArraySlice_l118_125 <= wReg);
  assign when_ArraySlice_l173_125 = (_zz_when_ArraySlice_l173_125_1 <= _zz_when_ArraySlice_l173_125_3);
  assign when_ArraySlice_l165_126 = (_zz_when_ArraySlice_l165_126 <= selectWriteFifo);
  assign when_ArraySlice_l166_126 = (_zz_when_ArraySlice_l166_126 <= _zz_when_ArraySlice_l166_126_2);
  assign _zz_when_ArraySlice_l112_126 = (wReg % _zz__zz_when_ArraySlice_l112_126);
  assign when_ArraySlice_l112_126 = (_zz_when_ArraySlice_l112_126 != 6'h0);
  assign when_ArraySlice_l113_126 = (7'h40 <= _zz_when_ArraySlice_l113_126);
  always @(*) begin
    if(when_ArraySlice_l112_126) begin
      if(when_ArraySlice_l113_126) begin
        _zz_when_ArraySlice_l173_126 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_126 = (_zz__zz_when_ArraySlice_l173_126 - _zz__zz_when_ArraySlice_l173_126_3);
      end
    end else begin
      if(when_ArraySlice_l118_126) begin
        _zz_when_ArraySlice_l173_126 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_126 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_126 = (_zz_when_ArraySlice_l118_126 <= wReg);
  assign when_ArraySlice_l173_126 = (_zz_when_ArraySlice_l173_126_1 <= _zz_when_ArraySlice_l173_126_3);
  assign when_ArraySlice_l165_127 = (_zz_when_ArraySlice_l165_127 <= selectWriteFifo);
  assign when_ArraySlice_l166_127 = (_zz_when_ArraySlice_l166_127 <= _zz_when_ArraySlice_l166_127_2);
  assign _zz_when_ArraySlice_l112_127 = (wReg % _zz__zz_when_ArraySlice_l112_127);
  assign when_ArraySlice_l112_127 = (_zz_when_ArraySlice_l112_127 != 6'h0);
  assign when_ArraySlice_l113_127 = (7'h40 <= _zz_when_ArraySlice_l113_127);
  always @(*) begin
    if(when_ArraySlice_l112_127) begin
      if(when_ArraySlice_l113_127) begin
        _zz_when_ArraySlice_l173_127 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_127 = (_zz__zz_when_ArraySlice_l173_127 - _zz__zz_when_ArraySlice_l173_127_3);
      end
    end else begin
      if(when_ArraySlice_l118_127) begin
        _zz_when_ArraySlice_l173_127 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_127 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_127 = (_zz_when_ArraySlice_l118_127 <= wReg);
  assign when_ArraySlice_l173_127 = (_zz_when_ArraySlice_l173_127_1 <= _zz_when_ArraySlice_l173_127_3);
  assign when_ArraySlice_l444_4 = (! ((((((_zz_when_ArraySlice_l444_4_1 && _zz_when_ArraySlice_l444_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l444_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l444_4_4 && _zz_when_ArraySlice_l444_4_5) && (debug_4_15 == _zz_when_ArraySlice_l444_4_6)) && (debug_5_15 == 1'b1)) && (debug_6_15 == 1'b1)) && (debug_7_15 == 1'b1))));
  assign outputStreamArrayData_4_fire_5 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l448_4 = ((_zz_when_ArraySlice_l448_4 == 13'h0) && outputStreamArrayData_4_fire_5);
  assign when_ArraySlice_l434_4 = (allowPadding_4 && (wReg <= _zz_when_ArraySlice_l434_4));
  assign outputStreamArrayData_4_fire_6 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l455_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l455_4_1);
  assign when_ArraySlice_l373_5 = (_zz_when_ArraySlice_l373_5 < wReg);
  assign when_ArraySlice_l374_5 = ((! holdReadOp_5) && (_zz_when_ArraySlice_l374_5 != 7'h0));
  assign _zz_outputStreamArrayData_5_valid = (selectReadFifo_5 + _zz__zz_outputStreamArrayData_5_valid);
  assign _zz_8 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_5_valid);
  assign _zz_io_pop_ready_5 = outputStreamArrayData_5_ready;
  assign when_ArraySlice_l379_5 = (! holdReadOp_5);
  assign outputStreamArrayData_5_fire = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l380_5 = ((_zz_when_ArraySlice_l380_5_1 < _zz_when_ArraySlice_l380_5_3) && outputStreamArrayData_5_fire);
  assign when_ArraySlice_l381_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l381_5);
  assign when_ArraySlice_l384_5 = (_zz_when_ArraySlice_l384_5 == 13'h0);
  assign outputStreamArrayData_5_fire_1 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l389_5 = ((_zz_when_ArraySlice_l389_5_1 == _zz_when_ArraySlice_l389_5_4) && outputStreamArrayData_5_fire_1);
  assign when_ArraySlice_l390_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l390_5);
  assign _zz_when_ArraySlice_l94_15 = (hReg % _zz__zz_when_ArraySlice_l94_15);
  assign when_ArraySlice_l94_15 = (_zz_when_ArraySlice_l94_15 != 6'h0);
  assign when_ArraySlice_l95_15 = (7'h40 <= _zz_when_ArraySlice_l95_15);
  always @(*) begin
    if(when_ArraySlice_l94_15) begin
      if(when_ArraySlice_l95_15) begin
        _zz_when_ArraySlice_l392_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_5 = (_zz__zz_when_ArraySlice_l392_5 - _zz__zz_when_ArraySlice_l392_5_3);
      end
    end else begin
      if(when_ArraySlice_l99_15) begin
        _zz_when_ArraySlice_l392_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_5 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_15 = (_zz_when_ArraySlice_l99_15 <= hReg);
  assign when_ArraySlice_l392_5 = (_zz_when_ArraySlice_l392_5_1 < _zz_when_ArraySlice_l392_5_4);
  always @(*) begin
    debug_0_16 = 1'b0;
    if(when_ArraySlice_l165_128) begin
      if(when_ArraySlice_l166_128) begin
        debug_0_16 = 1'b1;
      end else begin
        debug_0_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_128) begin
        debug_0_16 = 1'b1;
      end else begin
        debug_0_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_16 = 1'b0;
    if(when_ArraySlice_l165_129) begin
      if(when_ArraySlice_l166_129) begin
        debug_1_16 = 1'b1;
      end else begin
        debug_1_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_129) begin
        debug_1_16 = 1'b1;
      end else begin
        debug_1_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_16 = 1'b0;
    if(when_ArraySlice_l165_130) begin
      if(when_ArraySlice_l166_130) begin
        debug_2_16 = 1'b1;
      end else begin
        debug_2_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_130) begin
        debug_2_16 = 1'b1;
      end else begin
        debug_2_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_16 = 1'b0;
    if(when_ArraySlice_l165_131) begin
      if(when_ArraySlice_l166_131) begin
        debug_3_16 = 1'b1;
      end else begin
        debug_3_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_131) begin
        debug_3_16 = 1'b1;
      end else begin
        debug_3_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_16 = 1'b0;
    if(when_ArraySlice_l165_132) begin
      if(when_ArraySlice_l166_132) begin
        debug_4_16 = 1'b1;
      end else begin
        debug_4_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_132) begin
        debug_4_16 = 1'b1;
      end else begin
        debug_4_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_16 = 1'b0;
    if(when_ArraySlice_l165_133) begin
      if(when_ArraySlice_l166_133) begin
        debug_5_16 = 1'b1;
      end else begin
        debug_5_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_133) begin
        debug_5_16 = 1'b1;
      end else begin
        debug_5_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_16 = 1'b0;
    if(when_ArraySlice_l165_134) begin
      if(when_ArraySlice_l166_134) begin
        debug_6_16 = 1'b1;
      end else begin
        debug_6_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_134) begin
        debug_6_16 = 1'b1;
      end else begin
        debug_6_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_16 = 1'b0;
    if(when_ArraySlice_l165_135) begin
      if(when_ArraySlice_l166_135) begin
        debug_7_16 = 1'b1;
      end else begin
        debug_7_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_135) begin
        debug_7_16 = 1'b1;
      end else begin
        debug_7_16 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_128 = (_zz_when_ArraySlice_l165_128 <= selectWriteFifo);
  assign when_ArraySlice_l166_128 = (_zz_when_ArraySlice_l166_128 <= _zz_when_ArraySlice_l166_128_1);
  assign _zz_when_ArraySlice_l112_128 = (wReg % _zz__zz_when_ArraySlice_l112_128);
  assign when_ArraySlice_l112_128 = (_zz_when_ArraySlice_l112_128 != 6'h0);
  assign when_ArraySlice_l113_128 = (7'h40 <= _zz_when_ArraySlice_l113_128);
  always @(*) begin
    if(when_ArraySlice_l112_128) begin
      if(when_ArraySlice_l113_128) begin
        _zz_when_ArraySlice_l173_128 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_128 = (_zz__zz_when_ArraySlice_l173_128 - _zz__zz_when_ArraySlice_l173_128_3);
      end
    end else begin
      if(when_ArraySlice_l118_128) begin
        _zz_when_ArraySlice_l173_128 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_128 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_128 = (_zz_when_ArraySlice_l118_128 <= wReg);
  assign when_ArraySlice_l173_128 = (_zz_when_ArraySlice_l173_128_1 <= _zz_when_ArraySlice_l173_128_2);
  assign when_ArraySlice_l165_129 = (_zz_when_ArraySlice_l165_129 <= selectWriteFifo);
  assign when_ArraySlice_l166_129 = (_zz_when_ArraySlice_l166_129 <= _zz_when_ArraySlice_l166_129_1);
  assign _zz_when_ArraySlice_l112_129 = (wReg % _zz__zz_when_ArraySlice_l112_129);
  assign when_ArraySlice_l112_129 = (_zz_when_ArraySlice_l112_129 != 6'h0);
  assign when_ArraySlice_l113_129 = (7'h40 <= _zz_when_ArraySlice_l113_129);
  always @(*) begin
    if(when_ArraySlice_l112_129) begin
      if(when_ArraySlice_l113_129) begin
        _zz_when_ArraySlice_l173_129 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_129 = (_zz__zz_when_ArraySlice_l173_129 - _zz__zz_when_ArraySlice_l173_129_3);
      end
    end else begin
      if(when_ArraySlice_l118_129) begin
        _zz_when_ArraySlice_l173_129 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_129 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_129 = (_zz_when_ArraySlice_l118_129 <= wReg);
  assign when_ArraySlice_l173_129 = (_zz_when_ArraySlice_l173_129_1 <= _zz_when_ArraySlice_l173_129_3);
  assign when_ArraySlice_l165_130 = (_zz_when_ArraySlice_l165_130 <= selectWriteFifo);
  assign when_ArraySlice_l166_130 = (_zz_when_ArraySlice_l166_130 <= _zz_when_ArraySlice_l166_130_1);
  assign _zz_when_ArraySlice_l112_130 = (wReg % _zz__zz_when_ArraySlice_l112_130);
  assign when_ArraySlice_l112_130 = (_zz_when_ArraySlice_l112_130 != 6'h0);
  assign when_ArraySlice_l113_130 = (7'h40 <= _zz_when_ArraySlice_l113_130);
  always @(*) begin
    if(when_ArraySlice_l112_130) begin
      if(when_ArraySlice_l113_130) begin
        _zz_when_ArraySlice_l173_130 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_130 = (_zz__zz_when_ArraySlice_l173_130 - _zz__zz_when_ArraySlice_l173_130_3);
      end
    end else begin
      if(when_ArraySlice_l118_130) begin
        _zz_when_ArraySlice_l173_130 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_130 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_130 = (_zz_when_ArraySlice_l118_130 <= wReg);
  assign when_ArraySlice_l173_130 = (_zz_when_ArraySlice_l173_130_1 <= _zz_when_ArraySlice_l173_130_3);
  assign when_ArraySlice_l165_131 = (_zz_when_ArraySlice_l165_131 <= selectWriteFifo);
  assign when_ArraySlice_l166_131 = (_zz_when_ArraySlice_l166_131 <= _zz_when_ArraySlice_l166_131_1);
  assign _zz_when_ArraySlice_l112_131 = (wReg % _zz__zz_when_ArraySlice_l112_131);
  assign when_ArraySlice_l112_131 = (_zz_when_ArraySlice_l112_131 != 6'h0);
  assign when_ArraySlice_l113_131 = (7'h40 <= _zz_when_ArraySlice_l113_131);
  always @(*) begin
    if(when_ArraySlice_l112_131) begin
      if(when_ArraySlice_l113_131) begin
        _zz_when_ArraySlice_l173_131 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_131 = (_zz__zz_when_ArraySlice_l173_131 - _zz__zz_when_ArraySlice_l173_131_3);
      end
    end else begin
      if(when_ArraySlice_l118_131) begin
        _zz_when_ArraySlice_l173_131 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_131 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_131 = (_zz_when_ArraySlice_l118_131 <= wReg);
  assign when_ArraySlice_l173_131 = (_zz_when_ArraySlice_l173_131_1 <= _zz_when_ArraySlice_l173_131_3);
  assign when_ArraySlice_l165_132 = (_zz_when_ArraySlice_l165_132 <= selectWriteFifo);
  assign when_ArraySlice_l166_132 = (_zz_when_ArraySlice_l166_132 <= _zz_when_ArraySlice_l166_132_1);
  assign _zz_when_ArraySlice_l112_132 = (wReg % _zz__zz_when_ArraySlice_l112_132);
  assign when_ArraySlice_l112_132 = (_zz_when_ArraySlice_l112_132 != 6'h0);
  assign when_ArraySlice_l113_132 = (7'h40 <= _zz_when_ArraySlice_l113_132);
  always @(*) begin
    if(when_ArraySlice_l112_132) begin
      if(when_ArraySlice_l113_132) begin
        _zz_when_ArraySlice_l173_132 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_132 = (_zz__zz_when_ArraySlice_l173_132 - _zz__zz_when_ArraySlice_l173_132_3);
      end
    end else begin
      if(when_ArraySlice_l118_132) begin
        _zz_when_ArraySlice_l173_132 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_132 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_132 = (_zz_when_ArraySlice_l118_132 <= wReg);
  assign when_ArraySlice_l173_132 = (_zz_when_ArraySlice_l173_132_1 <= _zz_when_ArraySlice_l173_132_3);
  assign when_ArraySlice_l165_133 = (_zz_when_ArraySlice_l165_133 <= selectWriteFifo);
  assign when_ArraySlice_l166_133 = (_zz_when_ArraySlice_l166_133 <= _zz_when_ArraySlice_l166_133_2);
  assign _zz_when_ArraySlice_l112_133 = (wReg % _zz__zz_when_ArraySlice_l112_133);
  assign when_ArraySlice_l112_133 = (_zz_when_ArraySlice_l112_133 != 6'h0);
  assign when_ArraySlice_l113_133 = (7'h40 <= _zz_when_ArraySlice_l113_133);
  always @(*) begin
    if(when_ArraySlice_l112_133) begin
      if(when_ArraySlice_l113_133) begin
        _zz_when_ArraySlice_l173_133 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_133 = (_zz__zz_when_ArraySlice_l173_133 - _zz__zz_when_ArraySlice_l173_133_3);
      end
    end else begin
      if(when_ArraySlice_l118_133) begin
        _zz_when_ArraySlice_l173_133 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_133 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_133 = (_zz_when_ArraySlice_l118_133 <= wReg);
  assign when_ArraySlice_l173_133 = (_zz_when_ArraySlice_l173_133_1 <= _zz_when_ArraySlice_l173_133_3);
  assign when_ArraySlice_l165_134 = (_zz_when_ArraySlice_l165_134 <= selectWriteFifo);
  assign when_ArraySlice_l166_134 = (_zz_when_ArraySlice_l166_134 <= _zz_when_ArraySlice_l166_134_2);
  assign _zz_when_ArraySlice_l112_134 = (wReg % _zz__zz_when_ArraySlice_l112_134);
  assign when_ArraySlice_l112_134 = (_zz_when_ArraySlice_l112_134 != 6'h0);
  assign when_ArraySlice_l113_134 = (7'h40 <= _zz_when_ArraySlice_l113_134);
  always @(*) begin
    if(when_ArraySlice_l112_134) begin
      if(when_ArraySlice_l113_134) begin
        _zz_when_ArraySlice_l173_134 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_134 = (_zz__zz_when_ArraySlice_l173_134 - _zz__zz_when_ArraySlice_l173_134_3);
      end
    end else begin
      if(when_ArraySlice_l118_134) begin
        _zz_when_ArraySlice_l173_134 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_134 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_134 = (_zz_when_ArraySlice_l118_134 <= wReg);
  assign when_ArraySlice_l173_134 = (_zz_when_ArraySlice_l173_134_1 <= _zz_when_ArraySlice_l173_134_3);
  assign when_ArraySlice_l165_135 = (_zz_when_ArraySlice_l165_135 <= selectWriteFifo);
  assign when_ArraySlice_l166_135 = (_zz_when_ArraySlice_l166_135 <= _zz_when_ArraySlice_l166_135_2);
  assign _zz_when_ArraySlice_l112_135 = (wReg % _zz__zz_when_ArraySlice_l112_135);
  assign when_ArraySlice_l112_135 = (_zz_when_ArraySlice_l112_135 != 6'h0);
  assign when_ArraySlice_l113_135 = (7'h40 <= _zz_when_ArraySlice_l113_135);
  always @(*) begin
    if(when_ArraySlice_l112_135) begin
      if(when_ArraySlice_l113_135) begin
        _zz_when_ArraySlice_l173_135 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_135 = (_zz__zz_when_ArraySlice_l173_135 - _zz__zz_when_ArraySlice_l173_135_3);
      end
    end else begin
      if(when_ArraySlice_l118_135) begin
        _zz_when_ArraySlice_l173_135 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_135 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_135 = (_zz_when_ArraySlice_l118_135 <= wReg);
  assign when_ArraySlice_l173_135 = (_zz_when_ArraySlice_l173_135_1 <= _zz_when_ArraySlice_l173_135_3);
  assign when_ArraySlice_l398_5 = (! ((((((_zz_when_ArraySlice_l398_5_1 && _zz_when_ArraySlice_l398_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l398_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l398_5_4 && _zz_when_ArraySlice_l398_5_5) && (debug_4_16 == _zz_when_ArraySlice_l398_5_6)) && (debug_5_16 == 1'b1)) && (debug_6_16 == 1'b1)) && (debug_7_16 == 1'b1))));
  assign when_ArraySlice_l401_5 = (wReg <= _zz_when_ArraySlice_l401_5_1);
  assign when_ArraySlice_l405_5 = (_zz_when_ArraySlice_l405_5 == 13'h0);
  assign when_ArraySlice_l409_5 = (_zz_when_ArraySlice_l409_5 == 7'h0);
  assign outputStreamArrayData_5_fire_2 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l410_5 = ((handshakeTimes_5_value == _zz_when_ArraySlice_l410_5) && outputStreamArrayData_5_fire_2);
  assign _zz_when_ArraySlice_l94_16 = (hReg % _zz__zz_when_ArraySlice_l94_16);
  assign when_ArraySlice_l94_16 = (_zz_when_ArraySlice_l94_16 != 6'h0);
  assign when_ArraySlice_l95_16 = (7'h40 <= _zz_when_ArraySlice_l95_16);
  always @(*) begin
    if(when_ArraySlice_l94_16) begin
      if(when_ArraySlice_l95_16) begin
        _zz_when_ArraySlice_l412_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_5 = (_zz__zz_when_ArraySlice_l412_5 - _zz__zz_when_ArraySlice_l412_5_3);
      end
    end else begin
      if(when_ArraySlice_l99_16) begin
        _zz_when_ArraySlice_l412_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_5 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_16 = (_zz_when_ArraySlice_l99_16 <= hReg);
  assign when_ArraySlice_l412_5 = (_zz_when_ArraySlice_l412_5_1 < _zz_when_ArraySlice_l412_5_4);
  always @(*) begin
    debug_0_17 = 1'b0;
    if(when_ArraySlice_l165_136) begin
      if(when_ArraySlice_l166_136) begin
        debug_0_17 = 1'b1;
      end else begin
        debug_0_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_136) begin
        debug_0_17 = 1'b1;
      end else begin
        debug_0_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_17 = 1'b0;
    if(when_ArraySlice_l165_137) begin
      if(when_ArraySlice_l166_137) begin
        debug_1_17 = 1'b1;
      end else begin
        debug_1_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_137) begin
        debug_1_17 = 1'b1;
      end else begin
        debug_1_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_17 = 1'b0;
    if(when_ArraySlice_l165_138) begin
      if(when_ArraySlice_l166_138) begin
        debug_2_17 = 1'b1;
      end else begin
        debug_2_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_138) begin
        debug_2_17 = 1'b1;
      end else begin
        debug_2_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_17 = 1'b0;
    if(when_ArraySlice_l165_139) begin
      if(when_ArraySlice_l166_139) begin
        debug_3_17 = 1'b1;
      end else begin
        debug_3_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_139) begin
        debug_3_17 = 1'b1;
      end else begin
        debug_3_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_17 = 1'b0;
    if(when_ArraySlice_l165_140) begin
      if(when_ArraySlice_l166_140) begin
        debug_4_17 = 1'b1;
      end else begin
        debug_4_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_140) begin
        debug_4_17 = 1'b1;
      end else begin
        debug_4_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_17 = 1'b0;
    if(when_ArraySlice_l165_141) begin
      if(when_ArraySlice_l166_141) begin
        debug_5_17 = 1'b1;
      end else begin
        debug_5_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_141) begin
        debug_5_17 = 1'b1;
      end else begin
        debug_5_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_17 = 1'b0;
    if(when_ArraySlice_l165_142) begin
      if(when_ArraySlice_l166_142) begin
        debug_6_17 = 1'b1;
      end else begin
        debug_6_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_142) begin
        debug_6_17 = 1'b1;
      end else begin
        debug_6_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_17 = 1'b0;
    if(when_ArraySlice_l165_143) begin
      if(when_ArraySlice_l166_143) begin
        debug_7_17 = 1'b1;
      end else begin
        debug_7_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_143) begin
        debug_7_17 = 1'b1;
      end else begin
        debug_7_17 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_136 = (_zz_when_ArraySlice_l165_136 <= selectWriteFifo);
  assign when_ArraySlice_l166_136 = (_zz_when_ArraySlice_l166_136 <= _zz_when_ArraySlice_l166_136_1);
  assign _zz_when_ArraySlice_l112_136 = (wReg % _zz__zz_when_ArraySlice_l112_136);
  assign when_ArraySlice_l112_136 = (_zz_when_ArraySlice_l112_136 != 6'h0);
  assign when_ArraySlice_l113_136 = (7'h40 <= _zz_when_ArraySlice_l113_136);
  always @(*) begin
    if(when_ArraySlice_l112_136) begin
      if(when_ArraySlice_l113_136) begin
        _zz_when_ArraySlice_l173_136 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_136 = (_zz__zz_when_ArraySlice_l173_136 - _zz__zz_when_ArraySlice_l173_136_3);
      end
    end else begin
      if(when_ArraySlice_l118_136) begin
        _zz_when_ArraySlice_l173_136 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_136 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_136 = (_zz_when_ArraySlice_l118_136 <= wReg);
  assign when_ArraySlice_l173_136 = (_zz_when_ArraySlice_l173_136_1 <= _zz_when_ArraySlice_l173_136_2);
  assign when_ArraySlice_l165_137 = (_zz_when_ArraySlice_l165_137 <= selectWriteFifo);
  assign when_ArraySlice_l166_137 = (_zz_when_ArraySlice_l166_137 <= _zz_when_ArraySlice_l166_137_1);
  assign _zz_when_ArraySlice_l112_137 = (wReg % _zz__zz_when_ArraySlice_l112_137);
  assign when_ArraySlice_l112_137 = (_zz_when_ArraySlice_l112_137 != 6'h0);
  assign when_ArraySlice_l113_137 = (7'h40 <= _zz_when_ArraySlice_l113_137);
  always @(*) begin
    if(when_ArraySlice_l112_137) begin
      if(when_ArraySlice_l113_137) begin
        _zz_when_ArraySlice_l173_137 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_137 = (_zz__zz_when_ArraySlice_l173_137 - _zz__zz_when_ArraySlice_l173_137_3);
      end
    end else begin
      if(when_ArraySlice_l118_137) begin
        _zz_when_ArraySlice_l173_137 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_137 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_137 = (_zz_when_ArraySlice_l118_137 <= wReg);
  assign when_ArraySlice_l173_137 = (_zz_when_ArraySlice_l173_137_1 <= _zz_when_ArraySlice_l173_137_3);
  assign when_ArraySlice_l165_138 = (_zz_when_ArraySlice_l165_138 <= selectWriteFifo);
  assign when_ArraySlice_l166_138 = (_zz_when_ArraySlice_l166_138 <= _zz_when_ArraySlice_l166_138_1);
  assign _zz_when_ArraySlice_l112_138 = (wReg % _zz__zz_when_ArraySlice_l112_138);
  assign when_ArraySlice_l112_138 = (_zz_when_ArraySlice_l112_138 != 6'h0);
  assign when_ArraySlice_l113_138 = (7'h40 <= _zz_when_ArraySlice_l113_138);
  always @(*) begin
    if(when_ArraySlice_l112_138) begin
      if(when_ArraySlice_l113_138) begin
        _zz_when_ArraySlice_l173_138 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_138 = (_zz__zz_when_ArraySlice_l173_138 - _zz__zz_when_ArraySlice_l173_138_3);
      end
    end else begin
      if(when_ArraySlice_l118_138) begin
        _zz_when_ArraySlice_l173_138 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_138 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_138 = (_zz_when_ArraySlice_l118_138 <= wReg);
  assign when_ArraySlice_l173_138 = (_zz_when_ArraySlice_l173_138_1 <= _zz_when_ArraySlice_l173_138_3);
  assign when_ArraySlice_l165_139 = (_zz_when_ArraySlice_l165_139 <= selectWriteFifo);
  assign when_ArraySlice_l166_139 = (_zz_when_ArraySlice_l166_139 <= _zz_when_ArraySlice_l166_139_1);
  assign _zz_when_ArraySlice_l112_139 = (wReg % _zz__zz_when_ArraySlice_l112_139);
  assign when_ArraySlice_l112_139 = (_zz_when_ArraySlice_l112_139 != 6'h0);
  assign when_ArraySlice_l113_139 = (7'h40 <= _zz_when_ArraySlice_l113_139);
  always @(*) begin
    if(when_ArraySlice_l112_139) begin
      if(when_ArraySlice_l113_139) begin
        _zz_when_ArraySlice_l173_139 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_139 = (_zz__zz_when_ArraySlice_l173_139 - _zz__zz_when_ArraySlice_l173_139_3);
      end
    end else begin
      if(when_ArraySlice_l118_139) begin
        _zz_when_ArraySlice_l173_139 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_139 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_139 = (_zz_when_ArraySlice_l118_139 <= wReg);
  assign when_ArraySlice_l173_139 = (_zz_when_ArraySlice_l173_139_1 <= _zz_when_ArraySlice_l173_139_3);
  assign when_ArraySlice_l165_140 = (_zz_when_ArraySlice_l165_140 <= selectWriteFifo);
  assign when_ArraySlice_l166_140 = (_zz_when_ArraySlice_l166_140 <= _zz_when_ArraySlice_l166_140_1);
  assign _zz_when_ArraySlice_l112_140 = (wReg % _zz__zz_when_ArraySlice_l112_140);
  assign when_ArraySlice_l112_140 = (_zz_when_ArraySlice_l112_140 != 6'h0);
  assign when_ArraySlice_l113_140 = (7'h40 <= _zz_when_ArraySlice_l113_140);
  always @(*) begin
    if(when_ArraySlice_l112_140) begin
      if(when_ArraySlice_l113_140) begin
        _zz_when_ArraySlice_l173_140 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_140 = (_zz__zz_when_ArraySlice_l173_140 - _zz__zz_when_ArraySlice_l173_140_3);
      end
    end else begin
      if(when_ArraySlice_l118_140) begin
        _zz_when_ArraySlice_l173_140 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_140 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_140 = (_zz_when_ArraySlice_l118_140 <= wReg);
  assign when_ArraySlice_l173_140 = (_zz_when_ArraySlice_l173_140_1 <= _zz_when_ArraySlice_l173_140_3);
  assign when_ArraySlice_l165_141 = (_zz_when_ArraySlice_l165_141 <= selectWriteFifo);
  assign when_ArraySlice_l166_141 = (_zz_when_ArraySlice_l166_141 <= _zz_when_ArraySlice_l166_141_2);
  assign _zz_when_ArraySlice_l112_141 = (wReg % _zz__zz_when_ArraySlice_l112_141);
  assign when_ArraySlice_l112_141 = (_zz_when_ArraySlice_l112_141 != 6'h0);
  assign when_ArraySlice_l113_141 = (7'h40 <= _zz_when_ArraySlice_l113_141);
  always @(*) begin
    if(when_ArraySlice_l112_141) begin
      if(when_ArraySlice_l113_141) begin
        _zz_when_ArraySlice_l173_141 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_141 = (_zz__zz_when_ArraySlice_l173_141 - _zz__zz_when_ArraySlice_l173_141_3);
      end
    end else begin
      if(when_ArraySlice_l118_141) begin
        _zz_when_ArraySlice_l173_141 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_141 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_141 = (_zz_when_ArraySlice_l118_141 <= wReg);
  assign when_ArraySlice_l173_141 = (_zz_when_ArraySlice_l173_141_1 <= _zz_when_ArraySlice_l173_141_3);
  assign when_ArraySlice_l165_142 = (_zz_when_ArraySlice_l165_142 <= selectWriteFifo);
  assign when_ArraySlice_l166_142 = (_zz_when_ArraySlice_l166_142 <= _zz_when_ArraySlice_l166_142_2);
  assign _zz_when_ArraySlice_l112_142 = (wReg % _zz__zz_when_ArraySlice_l112_142);
  assign when_ArraySlice_l112_142 = (_zz_when_ArraySlice_l112_142 != 6'h0);
  assign when_ArraySlice_l113_142 = (7'h40 <= _zz_when_ArraySlice_l113_142);
  always @(*) begin
    if(when_ArraySlice_l112_142) begin
      if(when_ArraySlice_l113_142) begin
        _zz_when_ArraySlice_l173_142 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_142 = (_zz__zz_when_ArraySlice_l173_142 - _zz__zz_when_ArraySlice_l173_142_3);
      end
    end else begin
      if(when_ArraySlice_l118_142) begin
        _zz_when_ArraySlice_l173_142 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_142 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_142 = (_zz_when_ArraySlice_l118_142 <= wReg);
  assign when_ArraySlice_l173_142 = (_zz_when_ArraySlice_l173_142_1 <= _zz_when_ArraySlice_l173_142_3);
  assign when_ArraySlice_l165_143 = (_zz_when_ArraySlice_l165_143 <= selectWriteFifo);
  assign when_ArraySlice_l166_143 = (_zz_when_ArraySlice_l166_143 <= _zz_when_ArraySlice_l166_143_2);
  assign _zz_when_ArraySlice_l112_143 = (wReg % _zz__zz_when_ArraySlice_l112_143);
  assign when_ArraySlice_l112_143 = (_zz_when_ArraySlice_l112_143 != 6'h0);
  assign when_ArraySlice_l113_143 = (7'h40 <= _zz_when_ArraySlice_l113_143);
  always @(*) begin
    if(when_ArraySlice_l112_143) begin
      if(when_ArraySlice_l113_143) begin
        _zz_when_ArraySlice_l173_143 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_143 = (_zz__zz_when_ArraySlice_l173_143 - _zz__zz_when_ArraySlice_l173_143_3);
      end
    end else begin
      if(when_ArraySlice_l118_143) begin
        _zz_when_ArraySlice_l173_143 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_143 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_143 = (_zz_when_ArraySlice_l118_143 <= wReg);
  assign when_ArraySlice_l173_143 = (_zz_when_ArraySlice_l173_143_1 <= _zz_when_ArraySlice_l173_143_3);
  assign when_ArraySlice_l418_5 = (! ((((((_zz_when_ArraySlice_l418_5_1 && _zz_when_ArraySlice_l418_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l418_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l418_5_4 && _zz_when_ArraySlice_l418_5_5) && (debug_4_17 == _zz_when_ArraySlice_l418_5_6)) && (debug_5_17 == 1'b1)) && (debug_6_17 == 1'b1)) && (debug_7_17 == 1'b1))));
  assign when_ArraySlice_l421_5 = (wReg <= _zz_when_ArraySlice_l421_5_1);
  assign outputStreamArrayData_5_fire_3 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l425_5 = ((_zz_when_ArraySlice_l425_5 == 13'h0) && outputStreamArrayData_5_fire_3);
  assign outputStreamArrayData_5_fire_4 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l436_5 = ((handshakeTimes_5_value == _zz_when_ArraySlice_l436_5) && outputStreamArrayData_5_fire_4);
  assign _zz_when_ArraySlice_l94_17 = (hReg % _zz__zz_when_ArraySlice_l94_17);
  assign when_ArraySlice_l94_17 = (_zz_when_ArraySlice_l94_17 != 6'h0);
  assign when_ArraySlice_l95_17 = (7'h40 <= _zz_when_ArraySlice_l95_17);
  always @(*) begin
    if(when_ArraySlice_l94_17) begin
      if(when_ArraySlice_l95_17) begin
        _zz_when_ArraySlice_l437_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_5 = (_zz__zz_when_ArraySlice_l437_5 - _zz__zz_when_ArraySlice_l437_5_3);
      end
    end else begin
      if(when_ArraySlice_l99_17) begin
        _zz_when_ArraySlice_l437_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_5 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_17 = (_zz_when_ArraySlice_l99_17 <= hReg);
  assign when_ArraySlice_l437_5 = (_zz_when_ArraySlice_l437_5_1 < _zz_when_ArraySlice_l437_5_4);
  always @(*) begin
    debug_0_18 = 1'b0;
    if(when_ArraySlice_l165_144) begin
      if(when_ArraySlice_l166_144) begin
        debug_0_18 = 1'b1;
      end else begin
        debug_0_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_144) begin
        debug_0_18 = 1'b1;
      end else begin
        debug_0_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_18 = 1'b0;
    if(when_ArraySlice_l165_145) begin
      if(when_ArraySlice_l166_145) begin
        debug_1_18 = 1'b1;
      end else begin
        debug_1_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_145) begin
        debug_1_18 = 1'b1;
      end else begin
        debug_1_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_18 = 1'b0;
    if(when_ArraySlice_l165_146) begin
      if(when_ArraySlice_l166_146) begin
        debug_2_18 = 1'b1;
      end else begin
        debug_2_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_146) begin
        debug_2_18 = 1'b1;
      end else begin
        debug_2_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_18 = 1'b0;
    if(when_ArraySlice_l165_147) begin
      if(when_ArraySlice_l166_147) begin
        debug_3_18 = 1'b1;
      end else begin
        debug_3_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_147) begin
        debug_3_18 = 1'b1;
      end else begin
        debug_3_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_18 = 1'b0;
    if(when_ArraySlice_l165_148) begin
      if(when_ArraySlice_l166_148) begin
        debug_4_18 = 1'b1;
      end else begin
        debug_4_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_148) begin
        debug_4_18 = 1'b1;
      end else begin
        debug_4_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_18 = 1'b0;
    if(when_ArraySlice_l165_149) begin
      if(when_ArraySlice_l166_149) begin
        debug_5_18 = 1'b1;
      end else begin
        debug_5_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_149) begin
        debug_5_18 = 1'b1;
      end else begin
        debug_5_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_18 = 1'b0;
    if(when_ArraySlice_l165_150) begin
      if(when_ArraySlice_l166_150) begin
        debug_6_18 = 1'b1;
      end else begin
        debug_6_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_150) begin
        debug_6_18 = 1'b1;
      end else begin
        debug_6_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_18 = 1'b0;
    if(when_ArraySlice_l165_151) begin
      if(when_ArraySlice_l166_151) begin
        debug_7_18 = 1'b1;
      end else begin
        debug_7_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_151) begin
        debug_7_18 = 1'b1;
      end else begin
        debug_7_18 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_144 = (_zz_when_ArraySlice_l165_144 <= selectWriteFifo);
  assign when_ArraySlice_l166_144 = (_zz_when_ArraySlice_l166_144 <= _zz_when_ArraySlice_l166_144_1);
  assign _zz_when_ArraySlice_l112_144 = (wReg % _zz__zz_when_ArraySlice_l112_144);
  assign when_ArraySlice_l112_144 = (_zz_when_ArraySlice_l112_144 != 6'h0);
  assign when_ArraySlice_l113_144 = (7'h40 <= _zz_when_ArraySlice_l113_144);
  always @(*) begin
    if(when_ArraySlice_l112_144) begin
      if(when_ArraySlice_l113_144) begin
        _zz_when_ArraySlice_l173_144 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_144 = (_zz__zz_when_ArraySlice_l173_144 - _zz__zz_when_ArraySlice_l173_144_3);
      end
    end else begin
      if(when_ArraySlice_l118_144) begin
        _zz_when_ArraySlice_l173_144 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_144 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_144 = (_zz_when_ArraySlice_l118_144 <= wReg);
  assign when_ArraySlice_l173_144 = (_zz_when_ArraySlice_l173_144_1 <= _zz_when_ArraySlice_l173_144_2);
  assign when_ArraySlice_l165_145 = (_zz_when_ArraySlice_l165_145 <= selectWriteFifo);
  assign when_ArraySlice_l166_145 = (_zz_when_ArraySlice_l166_145 <= _zz_when_ArraySlice_l166_145_1);
  assign _zz_when_ArraySlice_l112_145 = (wReg % _zz__zz_when_ArraySlice_l112_145);
  assign when_ArraySlice_l112_145 = (_zz_when_ArraySlice_l112_145 != 6'h0);
  assign when_ArraySlice_l113_145 = (7'h40 <= _zz_when_ArraySlice_l113_145);
  always @(*) begin
    if(when_ArraySlice_l112_145) begin
      if(when_ArraySlice_l113_145) begin
        _zz_when_ArraySlice_l173_145 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_145 = (_zz__zz_when_ArraySlice_l173_145 - _zz__zz_when_ArraySlice_l173_145_3);
      end
    end else begin
      if(when_ArraySlice_l118_145) begin
        _zz_when_ArraySlice_l173_145 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_145 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_145 = (_zz_when_ArraySlice_l118_145 <= wReg);
  assign when_ArraySlice_l173_145 = (_zz_when_ArraySlice_l173_145_1 <= _zz_when_ArraySlice_l173_145_3);
  assign when_ArraySlice_l165_146 = (_zz_when_ArraySlice_l165_146 <= selectWriteFifo);
  assign when_ArraySlice_l166_146 = (_zz_when_ArraySlice_l166_146 <= _zz_when_ArraySlice_l166_146_1);
  assign _zz_when_ArraySlice_l112_146 = (wReg % _zz__zz_when_ArraySlice_l112_146);
  assign when_ArraySlice_l112_146 = (_zz_when_ArraySlice_l112_146 != 6'h0);
  assign when_ArraySlice_l113_146 = (7'h40 <= _zz_when_ArraySlice_l113_146);
  always @(*) begin
    if(when_ArraySlice_l112_146) begin
      if(when_ArraySlice_l113_146) begin
        _zz_when_ArraySlice_l173_146 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_146 = (_zz__zz_when_ArraySlice_l173_146 - _zz__zz_when_ArraySlice_l173_146_3);
      end
    end else begin
      if(when_ArraySlice_l118_146) begin
        _zz_when_ArraySlice_l173_146 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_146 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_146 = (_zz_when_ArraySlice_l118_146 <= wReg);
  assign when_ArraySlice_l173_146 = (_zz_when_ArraySlice_l173_146_1 <= _zz_when_ArraySlice_l173_146_3);
  assign when_ArraySlice_l165_147 = (_zz_when_ArraySlice_l165_147 <= selectWriteFifo);
  assign when_ArraySlice_l166_147 = (_zz_when_ArraySlice_l166_147 <= _zz_when_ArraySlice_l166_147_1);
  assign _zz_when_ArraySlice_l112_147 = (wReg % _zz__zz_when_ArraySlice_l112_147);
  assign when_ArraySlice_l112_147 = (_zz_when_ArraySlice_l112_147 != 6'h0);
  assign when_ArraySlice_l113_147 = (7'h40 <= _zz_when_ArraySlice_l113_147);
  always @(*) begin
    if(when_ArraySlice_l112_147) begin
      if(when_ArraySlice_l113_147) begin
        _zz_when_ArraySlice_l173_147 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_147 = (_zz__zz_when_ArraySlice_l173_147 - _zz__zz_when_ArraySlice_l173_147_3);
      end
    end else begin
      if(when_ArraySlice_l118_147) begin
        _zz_when_ArraySlice_l173_147 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_147 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_147 = (_zz_when_ArraySlice_l118_147 <= wReg);
  assign when_ArraySlice_l173_147 = (_zz_when_ArraySlice_l173_147_1 <= _zz_when_ArraySlice_l173_147_3);
  assign when_ArraySlice_l165_148 = (_zz_when_ArraySlice_l165_148 <= selectWriteFifo);
  assign when_ArraySlice_l166_148 = (_zz_when_ArraySlice_l166_148 <= _zz_when_ArraySlice_l166_148_1);
  assign _zz_when_ArraySlice_l112_148 = (wReg % _zz__zz_when_ArraySlice_l112_148);
  assign when_ArraySlice_l112_148 = (_zz_when_ArraySlice_l112_148 != 6'h0);
  assign when_ArraySlice_l113_148 = (7'h40 <= _zz_when_ArraySlice_l113_148);
  always @(*) begin
    if(when_ArraySlice_l112_148) begin
      if(when_ArraySlice_l113_148) begin
        _zz_when_ArraySlice_l173_148 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_148 = (_zz__zz_when_ArraySlice_l173_148 - _zz__zz_when_ArraySlice_l173_148_3);
      end
    end else begin
      if(when_ArraySlice_l118_148) begin
        _zz_when_ArraySlice_l173_148 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_148 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_148 = (_zz_when_ArraySlice_l118_148 <= wReg);
  assign when_ArraySlice_l173_148 = (_zz_when_ArraySlice_l173_148_1 <= _zz_when_ArraySlice_l173_148_3);
  assign when_ArraySlice_l165_149 = (_zz_when_ArraySlice_l165_149 <= selectWriteFifo);
  assign when_ArraySlice_l166_149 = (_zz_when_ArraySlice_l166_149 <= _zz_when_ArraySlice_l166_149_2);
  assign _zz_when_ArraySlice_l112_149 = (wReg % _zz__zz_when_ArraySlice_l112_149);
  assign when_ArraySlice_l112_149 = (_zz_when_ArraySlice_l112_149 != 6'h0);
  assign when_ArraySlice_l113_149 = (7'h40 <= _zz_when_ArraySlice_l113_149);
  always @(*) begin
    if(when_ArraySlice_l112_149) begin
      if(when_ArraySlice_l113_149) begin
        _zz_when_ArraySlice_l173_149 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_149 = (_zz__zz_when_ArraySlice_l173_149 - _zz__zz_when_ArraySlice_l173_149_3);
      end
    end else begin
      if(when_ArraySlice_l118_149) begin
        _zz_when_ArraySlice_l173_149 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_149 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_149 = (_zz_when_ArraySlice_l118_149 <= wReg);
  assign when_ArraySlice_l173_149 = (_zz_when_ArraySlice_l173_149_1 <= _zz_when_ArraySlice_l173_149_3);
  assign when_ArraySlice_l165_150 = (_zz_when_ArraySlice_l165_150 <= selectWriteFifo);
  assign when_ArraySlice_l166_150 = (_zz_when_ArraySlice_l166_150 <= _zz_when_ArraySlice_l166_150_2);
  assign _zz_when_ArraySlice_l112_150 = (wReg % _zz__zz_when_ArraySlice_l112_150);
  assign when_ArraySlice_l112_150 = (_zz_when_ArraySlice_l112_150 != 6'h0);
  assign when_ArraySlice_l113_150 = (7'h40 <= _zz_when_ArraySlice_l113_150);
  always @(*) begin
    if(when_ArraySlice_l112_150) begin
      if(when_ArraySlice_l113_150) begin
        _zz_when_ArraySlice_l173_150 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_150 = (_zz__zz_when_ArraySlice_l173_150 - _zz__zz_when_ArraySlice_l173_150_3);
      end
    end else begin
      if(when_ArraySlice_l118_150) begin
        _zz_when_ArraySlice_l173_150 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_150 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_150 = (_zz_when_ArraySlice_l118_150 <= wReg);
  assign when_ArraySlice_l173_150 = (_zz_when_ArraySlice_l173_150_1 <= _zz_when_ArraySlice_l173_150_3);
  assign when_ArraySlice_l165_151 = (_zz_when_ArraySlice_l165_151 <= selectWriteFifo);
  assign when_ArraySlice_l166_151 = (_zz_when_ArraySlice_l166_151 <= _zz_when_ArraySlice_l166_151_2);
  assign _zz_when_ArraySlice_l112_151 = (wReg % _zz__zz_when_ArraySlice_l112_151);
  assign when_ArraySlice_l112_151 = (_zz_when_ArraySlice_l112_151 != 6'h0);
  assign when_ArraySlice_l113_151 = (7'h40 <= _zz_when_ArraySlice_l113_151);
  always @(*) begin
    if(when_ArraySlice_l112_151) begin
      if(when_ArraySlice_l113_151) begin
        _zz_when_ArraySlice_l173_151 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_151 = (_zz__zz_when_ArraySlice_l173_151 - _zz__zz_when_ArraySlice_l173_151_3);
      end
    end else begin
      if(when_ArraySlice_l118_151) begin
        _zz_when_ArraySlice_l173_151 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_151 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_151 = (_zz_when_ArraySlice_l118_151 <= wReg);
  assign when_ArraySlice_l173_151 = (_zz_when_ArraySlice_l173_151_1 <= _zz_when_ArraySlice_l173_151_3);
  assign when_ArraySlice_l444_5 = (! ((((((_zz_when_ArraySlice_l444_5_1 && _zz_when_ArraySlice_l444_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l444_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l444_5_4 && _zz_when_ArraySlice_l444_5_5) && (debug_4_18 == _zz_when_ArraySlice_l444_5_6)) && (debug_5_18 == 1'b1)) && (debug_6_18 == 1'b1)) && (debug_7_18 == 1'b1))));
  assign outputStreamArrayData_5_fire_5 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l448_5 = ((_zz_when_ArraySlice_l448_5 == 13'h0) && outputStreamArrayData_5_fire_5);
  assign when_ArraySlice_l434_5 = (allowPadding_5 && (wReg <= _zz_when_ArraySlice_l434_5));
  assign outputStreamArrayData_5_fire_6 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l455_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l455_5);
  assign when_ArraySlice_l373_6 = (_zz_when_ArraySlice_l373_6 < wReg);
  assign when_ArraySlice_l374_6 = ((! holdReadOp_6) && (_zz_when_ArraySlice_l374_6 != 7'h0));
  assign _zz_outputStreamArrayData_6_valid = (selectReadFifo_6 + _zz__zz_outputStreamArrayData_6_valid);
  assign _zz_9 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_6_valid);
  assign _zz_io_pop_ready_6 = outputStreamArrayData_6_ready;
  assign when_ArraySlice_l379_6 = (! holdReadOp_6);
  assign outputStreamArrayData_6_fire = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l380_6 = ((_zz_when_ArraySlice_l380_6 < _zz_when_ArraySlice_l380_6_2) && outputStreamArrayData_6_fire);
  assign when_ArraySlice_l381_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l381_6);
  assign when_ArraySlice_l384_6 = (_zz_when_ArraySlice_l384_6 == 13'h0);
  assign outputStreamArrayData_6_fire_1 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l389_6 = ((_zz_when_ArraySlice_l389_6 == _zz_when_ArraySlice_l389_6_3) && outputStreamArrayData_6_fire_1);
  assign when_ArraySlice_l390_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l390_6);
  assign _zz_when_ArraySlice_l94_18 = (hReg % _zz__zz_when_ArraySlice_l94_18);
  assign when_ArraySlice_l94_18 = (_zz_when_ArraySlice_l94_18 != 6'h0);
  assign when_ArraySlice_l95_18 = (7'h40 <= _zz_when_ArraySlice_l95_18);
  always @(*) begin
    if(when_ArraySlice_l94_18) begin
      if(when_ArraySlice_l95_18) begin
        _zz_when_ArraySlice_l392_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_6 = (_zz__zz_when_ArraySlice_l392_6 - _zz__zz_when_ArraySlice_l392_6_3);
      end
    end else begin
      if(when_ArraySlice_l99_18) begin
        _zz_when_ArraySlice_l392_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_6 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_18 = (_zz_when_ArraySlice_l99_18 <= hReg);
  assign when_ArraySlice_l392_6 = (_zz_when_ArraySlice_l392_6_1 < _zz_when_ArraySlice_l392_6_4);
  always @(*) begin
    debug_0_19 = 1'b0;
    if(when_ArraySlice_l165_152) begin
      if(when_ArraySlice_l166_152) begin
        debug_0_19 = 1'b1;
      end else begin
        debug_0_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_152) begin
        debug_0_19 = 1'b1;
      end else begin
        debug_0_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_19 = 1'b0;
    if(when_ArraySlice_l165_153) begin
      if(when_ArraySlice_l166_153) begin
        debug_1_19 = 1'b1;
      end else begin
        debug_1_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_153) begin
        debug_1_19 = 1'b1;
      end else begin
        debug_1_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_19 = 1'b0;
    if(when_ArraySlice_l165_154) begin
      if(when_ArraySlice_l166_154) begin
        debug_2_19 = 1'b1;
      end else begin
        debug_2_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_154) begin
        debug_2_19 = 1'b1;
      end else begin
        debug_2_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_19 = 1'b0;
    if(when_ArraySlice_l165_155) begin
      if(when_ArraySlice_l166_155) begin
        debug_3_19 = 1'b1;
      end else begin
        debug_3_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_155) begin
        debug_3_19 = 1'b1;
      end else begin
        debug_3_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_19 = 1'b0;
    if(when_ArraySlice_l165_156) begin
      if(when_ArraySlice_l166_156) begin
        debug_4_19 = 1'b1;
      end else begin
        debug_4_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_156) begin
        debug_4_19 = 1'b1;
      end else begin
        debug_4_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_19 = 1'b0;
    if(when_ArraySlice_l165_157) begin
      if(when_ArraySlice_l166_157) begin
        debug_5_19 = 1'b1;
      end else begin
        debug_5_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_157) begin
        debug_5_19 = 1'b1;
      end else begin
        debug_5_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_19 = 1'b0;
    if(when_ArraySlice_l165_158) begin
      if(when_ArraySlice_l166_158) begin
        debug_6_19 = 1'b1;
      end else begin
        debug_6_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_158) begin
        debug_6_19 = 1'b1;
      end else begin
        debug_6_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_19 = 1'b0;
    if(when_ArraySlice_l165_159) begin
      if(when_ArraySlice_l166_159) begin
        debug_7_19 = 1'b1;
      end else begin
        debug_7_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_159) begin
        debug_7_19 = 1'b1;
      end else begin
        debug_7_19 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_152 = (_zz_when_ArraySlice_l165_152 <= selectWriteFifo);
  assign when_ArraySlice_l166_152 = (_zz_when_ArraySlice_l166_152 <= _zz_when_ArraySlice_l166_152_1);
  assign _zz_when_ArraySlice_l112_152 = (wReg % _zz__zz_when_ArraySlice_l112_152);
  assign when_ArraySlice_l112_152 = (_zz_when_ArraySlice_l112_152 != 6'h0);
  assign when_ArraySlice_l113_152 = (7'h40 <= _zz_when_ArraySlice_l113_152);
  always @(*) begin
    if(when_ArraySlice_l112_152) begin
      if(when_ArraySlice_l113_152) begin
        _zz_when_ArraySlice_l173_152 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_152 = (_zz__zz_when_ArraySlice_l173_152 - _zz__zz_when_ArraySlice_l173_152_3);
      end
    end else begin
      if(when_ArraySlice_l118_152) begin
        _zz_when_ArraySlice_l173_152 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_152 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_152 = (_zz_when_ArraySlice_l118_152 <= wReg);
  assign when_ArraySlice_l173_152 = (_zz_when_ArraySlice_l173_152_1 <= _zz_when_ArraySlice_l173_152_2);
  assign when_ArraySlice_l165_153 = (_zz_when_ArraySlice_l165_153 <= selectWriteFifo);
  assign when_ArraySlice_l166_153 = (_zz_when_ArraySlice_l166_153 <= _zz_when_ArraySlice_l166_153_1);
  assign _zz_when_ArraySlice_l112_153 = (wReg % _zz__zz_when_ArraySlice_l112_153);
  assign when_ArraySlice_l112_153 = (_zz_when_ArraySlice_l112_153 != 6'h0);
  assign when_ArraySlice_l113_153 = (7'h40 <= _zz_when_ArraySlice_l113_153);
  always @(*) begin
    if(when_ArraySlice_l112_153) begin
      if(when_ArraySlice_l113_153) begin
        _zz_when_ArraySlice_l173_153 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_153 = (_zz__zz_when_ArraySlice_l173_153 - _zz__zz_when_ArraySlice_l173_153_3);
      end
    end else begin
      if(when_ArraySlice_l118_153) begin
        _zz_when_ArraySlice_l173_153 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_153 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_153 = (_zz_when_ArraySlice_l118_153 <= wReg);
  assign when_ArraySlice_l173_153 = (_zz_when_ArraySlice_l173_153_1 <= _zz_when_ArraySlice_l173_153_3);
  assign when_ArraySlice_l165_154 = (_zz_when_ArraySlice_l165_154 <= selectWriteFifo);
  assign when_ArraySlice_l166_154 = (_zz_when_ArraySlice_l166_154 <= _zz_when_ArraySlice_l166_154_1);
  assign _zz_when_ArraySlice_l112_154 = (wReg % _zz__zz_when_ArraySlice_l112_154);
  assign when_ArraySlice_l112_154 = (_zz_when_ArraySlice_l112_154 != 6'h0);
  assign when_ArraySlice_l113_154 = (7'h40 <= _zz_when_ArraySlice_l113_154);
  always @(*) begin
    if(when_ArraySlice_l112_154) begin
      if(when_ArraySlice_l113_154) begin
        _zz_when_ArraySlice_l173_154 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_154 = (_zz__zz_when_ArraySlice_l173_154 - _zz__zz_when_ArraySlice_l173_154_3);
      end
    end else begin
      if(when_ArraySlice_l118_154) begin
        _zz_when_ArraySlice_l173_154 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_154 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_154 = (_zz_when_ArraySlice_l118_154 <= wReg);
  assign when_ArraySlice_l173_154 = (_zz_when_ArraySlice_l173_154_1 <= _zz_when_ArraySlice_l173_154_3);
  assign when_ArraySlice_l165_155 = (_zz_when_ArraySlice_l165_155 <= selectWriteFifo);
  assign when_ArraySlice_l166_155 = (_zz_when_ArraySlice_l166_155 <= _zz_when_ArraySlice_l166_155_1);
  assign _zz_when_ArraySlice_l112_155 = (wReg % _zz__zz_when_ArraySlice_l112_155);
  assign when_ArraySlice_l112_155 = (_zz_when_ArraySlice_l112_155 != 6'h0);
  assign when_ArraySlice_l113_155 = (7'h40 <= _zz_when_ArraySlice_l113_155);
  always @(*) begin
    if(when_ArraySlice_l112_155) begin
      if(when_ArraySlice_l113_155) begin
        _zz_when_ArraySlice_l173_155 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_155 = (_zz__zz_when_ArraySlice_l173_155 - _zz__zz_when_ArraySlice_l173_155_3);
      end
    end else begin
      if(when_ArraySlice_l118_155) begin
        _zz_when_ArraySlice_l173_155 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_155 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_155 = (_zz_when_ArraySlice_l118_155 <= wReg);
  assign when_ArraySlice_l173_155 = (_zz_when_ArraySlice_l173_155_1 <= _zz_when_ArraySlice_l173_155_3);
  assign when_ArraySlice_l165_156 = (_zz_when_ArraySlice_l165_156 <= selectWriteFifo);
  assign when_ArraySlice_l166_156 = (_zz_when_ArraySlice_l166_156 <= _zz_when_ArraySlice_l166_156_1);
  assign _zz_when_ArraySlice_l112_156 = (wReg % _zz__zz_when_ArraySlice_l112_156);
  assign when_ArraySlice_l112_156 = (_zz_when_ArraySlice_l112_156 != 6'h0);
  assign when_ArraySlice_l113_156 = (7'h40 <= _zz_when_ArraySlice_l113_156);
  always @(*) begin
    if(when_ArraySlice_l112_156) begin
      if(when_ArraySlice_l113_156) begin
        _zz_when_ArraySlice_l173_156 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_156 = (_zz__zz_when_ArraySlice_l173_156 - _zz__zz_when_ArraySlice_l173_156_3);
      end
    end else begin
      if(when_ArraySlice_l118_156) begin
        _zz_when_ArraySlice_l173_156 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_156 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_156 = (_zz_when_ArraySlice_l118_156 <= wReg);
  assign when_ArraySlice_l173_156 = (_zz_when_ArraySlice_l173_156_1 <= _zz_when_ArraySlice_l173_156_3);
  assign when_ArraySlice_l165_157 = (_zz_when_ArraySlice_l165_157 <= selectWriteFifo);
  assign when_ArraySlice_l166_157 = (_zz_when_ArraySlice_l166_157 <= _zz_when_ArraySlice_l166_157_2);
  assign _zz_when_ArraySlice_l112_157 = (wReg % _zz__zz_when_ArraySlice_l112_157);
  assign when_ArraySlice_l112_157 = (_zz_when_ArraySlice_l112_157 != 6'h0);
  assign when_ArraySlice_l113_157 = (7'h40 <= _zz_when_ArraySlice_l113_157);
  always @(*) begin
    if(when_ArraySlice_l112_157) begin
      if(when_ArraySlice_l113_157) begin
        _zz_when_ArraySlice_l173_157 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_157 = (_zz__zz_when_ArraySlice_l173_157 - _zz__zz_when_ArraySlice_l173_157_3);
      end
    end else begin
      if(when_ArraySlice_l118_157) begin
        _zz_when_ArraySlice_l173_157 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_157 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_157 = (_zz_when_ArraySlice_l118_157 <= wReg);
  assign when_ArraySlice_l173_157 = (_zz_when_ArraySlice_l173_157_1 <= _zz_when_ArraySlice_l173_157_3);
  assign when_ArraySlice_l165_158 = (_zz_when_ArraySlice_l165_158 <= selectWriteFifo);
  assign when_ArraySlice_l166_158 = (_zz_when_ArraySlice_l166_158 <= _zz_when_ArraySlice_l166_158_2);
  assign _zz_when_ArraySlice_l112_158 = (wReg % _zz__zz_when_ArraySlice_l112_158);
  assign when_ArraySlice_l112_158 = (_zz_when_ArraySlice_l112_158 != 6'h0);
  assign when_ArraySlice_l113_158 = (7'h40 <= _zz_when_ArraySlice_l113_158);
  always @(*) begin
    if(when_ArraySlice_l112_158) begin
      if(when_ArraySlice_l113_158) begin
        _zz_when_ArraySlice_l173_158 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_158 = (_zz__zz_when_ArraySlice_l173_158 - _zz__zz_when_ArraySlice_l173_158_3);
      end
    end else begin
      if(when_ArraySlice_l118_158) begin
        _zz_when_ArraySlice_l173_158 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_158 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_158 = (_zz_when_ArraySlice_l118_158 <= wReg);
  assign when_ArraySlice_l173_158 = (_zz_when_ArraySlice_l173_158_1 <= _zz_when_ArraySlice_l173_158_3);
  assign when_ArraySlice_l165_159 = (_zz_when_ArraySlice_l165_159 <= selectWriteFifo);
  assign when_ArraySlice_l166_159 = (_zz_when_ArraySlice_l166_159 <= _zz_when_ArraySlice_l166_159_2);
  assign _zz_when_ArraySlice_l112_159 = (wReg % _zz__zz_when_ArraySlice_l112_159);
  assign when_ArraySlice_l112_159 = (_zz_when_ArraySlice_l112_159 != 6'h0);
  assign when_ArraySlice_l113_159 = (7'h40 <= _zz_when_ArraySlice_l113_159);
  always @(*) begin
    if(when_ArraySlice_l112_159) begin
      if(when_ArraySlice_l113_159) begin
        _zz_when_ArraySlice_l173_159 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_159 = (_zz__zz_when_ArraySlice_l173_159 - _zz__zz_when_ArraySlice_l173_159_3);
      end
    end else begin
      if(when_ArraySlice_l118_159) begin
        _zz_when_ArraySlice_l173_159 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_159 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_159 = (_zz_when_ArraySlice_l118_159 <= wReg);
  assign when_ArraySlice_l173_159 = (_zz_when_ArraySlice_l173_159_1 <= _zz_when_ArraySlice_l173_159_3);
  assign when_ArraySlice_l398_6 = (! ((((((_zz_when_ArraySlice_l398_6_1 && _zz_when_ArraySlice_l398_6_2) && (holdReadOp_4 == _zz_when_ArraySlice_l398_6_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l398_6_4 && _zz_when_ArraySlice_l398_6_5) && (debug_4_19 == _zz_when_ArraySlice_l398_6_6)) && (debug_5_19 == 1'b1)) && (debug_6_19 == 1'b1)) && (debug_7_19 == 1'b1))));
  assign when_ArraySlice_l401_6 = (wReg <= _zz_when_ArraySlice_l401_6_1);
  assign when_ArraySlice_l405_6 = (_zz_when_ArraySlice_l405_6 == 13'h0);
  assign when_ArraySlice_l409_6 = (_zz_when_ArraySlice_l409_6 == 7'h0);
  assign outputStreamArrayData_6_fire_2 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l410_6 = ((handshakeTimes_6_value == _zz_when_ArraySlice_l410_6) && outputStreamArrayData_6_fire_2);
  assign _zz_when_ArraySlice_l94_19 = (hReg % _zz__zz_when_ArraySlice_l94_19);
  assign when_ArraySlice_l94_19 = (_zz_when_ArraySlice_l94_19 != 6'h0);
  assign when_ArraySlice_l95_19 = (7'h40 <= _zz_when_ArraySlice_l95_19);
  always @(*) begin
    if(when_ArraySlice_l94_19) begin
      if(when_ArraySlice_l95_19) begin
        _zz_when_ArraySlice_l412_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_6 = (_zz__zz_when_ArraySlice_l412_6 - _zz__zz_when_ArraySlice_l412_6_3);
      end
    end else begin
      if(when_ArraySlice_l99_19) begin
        _zz_when_ArraySlice_l412_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_6 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_19 = (_zz_when_ArraySlice_l99_19 <= hReg);
  assign when_ArraySlice_l412_6 = (_zz_when_ArraySlice_l412_6_1 < _zz_when_ArraySlice_l412_6_4);
  always @(*) begin
    debug_0_20 = 1'b0;
    if(when_ArraySlice_l165_160) begin
      if(when_ArraySlice_l166_160) begin
        debug_0_20 = 1'b1;
      end else begin
        debug_0_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_160) begin
        debug_0_20 = 1'b1;
      end else begin
        debug_0_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_20 = 1'b0;
    if(when_ArraySlice_l165_161) begin
      if(when_ArraySlice_l166_161) begin
        debug_1_20 = 1'b1;
      end else begin
        debug_1_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_161) begin
        debug_1_20 = 1'b1;
      end else begin
        debug_1_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_20 = 1'b0;
    if(when_ArraySlice_l165_162) begin
      if(when_ArraySlice_l166_162) begin
        debug_2_20 = 1'b1;
      end else begin
        debug_2_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_162) begin
        debug_2_20 = 1'b1;
      end else begin
        debug_2_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_20 = 1'b0;
    if(when_ArraySlice_l165_163) begin
      if(when_ArraySlice_l166_163) begin
        debug_3_20 = 1'b1;
      end else begin
        debug_3_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_163) begin
        debug_3_20 = 1'b1;
      end else begin
        debug_3_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_20 = 1'b0;
    if(when_ArraySlice_l165_164) begin
      if(when_ArraySlice_l166_164) begin
        debug_4_20 = 1'b1;
      end else begin
        debug_4_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_164) begin
        debug_4_20 = 1'b1;
      end else begin
        debug_4_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_20 = 1'b0;
    if(when_ArraySlice_l165_165) begin
      if(when_ArraySlice_l166_165) begin
        debug_5_20 = 1'b1;
      end else begin
        debug_5_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_165) begin
        debug_5_20 = 1'b1;
      end else begin
        debug_5_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_20 = 1'b0;
    if(when_ArraySlice_l165_166) begin
      if(when_ArraySlice_l166_166) begin
        debug_6_20 = 1'b1;
      end else begin
        debug_6_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_166) begin
        debug_6_20 = 1'b1;
      end else begin
        debug_6_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_20 = 1'b0;
    if(when_ArraySlice_l165_167) begin
      if(when_ArraySlice_l166_167) begin
        debug_7_20 = 1'b1;
      end else begin
        debug_7_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_167) begin
        debug_7_20 = 1'b1;
      end else begin
        debug_7_20 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_160 = (_zz_when_ArraySlice_l165_160 <= selectWriteFifo);
  assign when_ArraySlice_l166_160 = (_zz_when_ArraySlice_l166_160 <= _zz_when_ArraySlice_l166_160_1);
  assign _zz_when_ArraySlice_l112_160 = (wReg % _zz__zz_when_ArraySlice_l112_160);
  assign when_ArraySlice_l112_160 = (_zz_when_ArraySlice_l112_160 != 6'h0);
  assign when_ArraySlice_l113_160 = (7'h40 <= _zz_when_ArraySlice_l113_160);
  always @(*) begin
    if(when_ArraySlice_l112_160) begin
      if(when_ArraySlice_l113_160) begin
        _zz_when_ArraySlice_l173_160 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_160 = (_zz__zz_when_ArraySlice_l173_160 - _zz__zz_when_ArraySlice_l173_160_3);
      end
    end else begin
      if(when_ArraySlice_l118_160) begin
        _zz_when_ArraySlice_l173_160 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_160 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_160 = (_zz_when_ArraySlice_l118_160 <= wReg);
  assign when_ArraySlice_l173_160 = (_zz_when_ArraySlice_l173_160_1 <= _zz_when_ArraySlice_l173_160_2);
  assign when_ArraySlice_l165_161 = (_zz_when_ArraySlice_l165_161 <= selectWriteFifo);
  assign when_ArraySlice_l166_161 = (_zz_when_ArraySlice_l166_161 <= _zz_when_ArraySlice_l166_161_1);
  assign _zz_when_ArraySlice_l112_161 = (wReg % _zz__zz_when_ArraySlice_l112_161);
  assign when_ArraySlice_l112_161 = (_zz_when_ArraySlice_l112_161 != 6'h0);
  assign when_ArraySlice_l113_161 = (7'h40 <= _zz_when_ArraySlice_l113_161);
  always @(*) begin
    if(when_ArraySlice_l112_161) begin
      if(when_ArraySlice_l113_161) begin
        _zz_when_ArraySlice_l173_161 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_161 = (_zz__zz_when_ArraySlice_l173_161 - _zz__zz_when_ArraySlice_l173_161_3);
      end
    end else begin
      if(when_ArraySlice_l118_161) begin
        _zz_when_ArraySlice_l173_161 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_161 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_161 = (_zz_when_ArraySlice_l118_161 <= wReg);
  assign when_ArraySlice_l173_161 = (_zz_when_ArraySlice_l173_161_1 <= _zz_when_ArraySlice_l173_161_3);
  assign when_ArraySlice_l165_162 = (_zz_when_ArraySlice_l165_162 <= selectWriteFifo);
  assign when_ArraySlice_l166_162 = (_zz_when_ArraySlice_l166_162 <= _zz_when_ArraySlice_l166_162_1);
  assign _zz_when_ArraySlice_l112_162 = (wReg % _zz__zz_when_ArraySlice_l112_162);
  assign when_ArraySlice_l112_162 = (_zz_when_ArraySlice_l112_162 != 6'h0);
  assign when_ArraySlice_l113_162 = (7'h40 <= _zz_when_ArraySlice_l113_162);
  always @(*) begin
    if(when_ArraySlice_l112_162) begin
      if(when_ArraySlice_l113_162) begin
        _zz_when_ArraySlice_l173_162 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_162 = (_zz__zz_when_ArraySlice_l173_162 - _zz__zz_when_ArraySlice_l173_162_3);
      end
    end else begin
      if(when_ArraySlice_l118_162) begin
        _zz_when_ArraySlice_l173_162 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_162 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_162 = (_zz_when_ArraySlice_l118_162 <= wReg);
  assign when_ArraySlice_l173_162 = (_zz_when_ArraySlice_l173_162_1 <= _zz_when_ArraySlice_l173_162_3);
  assign when_ArraySlice_l165_163 = (_zz_when_ArraySlice_l165_163 <= selectWriteFifo);
  assign when_ArraySlice_l166_163 = (_zz_when_ArraySlice_l166_163 <= _zz_when_ArraySlice_l166_163_1);
  assign _zz_when_ArraySlice_l112_163 = (wReg % _zz__zz_when_ArraySlice_l112_163);
  assign when_ArraySlice_l112_163 = (_zz_when_ArraySlice_l112_163 != 6'h0);
  assign when_ArraySlice_l113_163 = (7'h40 <= _zz_when_ArraySlice_l113_163);
  always @(*) begin
    if(when_ArraySlice_l112_163) begin
      if(when_ArraySlice_l113_163) begin
        _zz_when_ArraySlice_l173_163 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_163 = (_zz__zz_when_ArraySlice_l173_163 - _zz__zz_when_ArraySlice_l173_163_3);
      end
    end else begin
      if(when_ArraySlice_l118_163) begin
        _zz_when_ArraySlice_l173_163 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_163 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_163 = (_zz_when_ArraySlice_l118_163 <= wReg);
  assign when_ArraySlice_l173_163 = (_zz_when_ArraySlice_l173_163_1 <= _zz_when_ArraySlice_l173_163_3);
  assign when_ArraySlice_l165_164 = (_zz_when_ArraySlice_l165_164 <= selectWriteFifo);
  assign when_ArraySlice_l166_164 = (_zz_when_ArraySlice_l166_164 <= _zz_when_ArraySlice_l166_164_1);
  assign _zz_when_ArraySlice_l112_164 = (wReg % _zz__zz_when_ArraySlice_l112_164);
  assign when_ArraySlice_l112_164 = (_zz_when_ArraySlice_l112_164 != 6'h0);
  assign when_ArraySlice_l113_164 = (7'h40 <= _zz_when_ArraySlice_l113_164);
  always @(*) begin
    if(when_ArraySlice_l112_164) begin
      if(when_ArraySlice_l113_164) begin
        _zz_when_ArraySlice_l173_164 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_164 = (_zz__zz_when_ArraySlice_l173_164 - _zz__zz_when_ArraySlice_l173_164_3);
      end
    end else begin
      if(when_ArraySlice_l118_164) begin
        _zz_when_ArraySlice_l173_164 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_164 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_164 = (_zz_when_ArraySlice_l118_164 <= wReg);
  assign when_ArraySlice_l173_164 = (_zz_when_ArraySlice_l173_164_1 <= _zz_when_ArraySlice_l173_164_3);
  assign when_ArraySlice_l165_165 = (_zz_when_ArraySlice_l165_165 <= selectWriteFifo);
  assign when_ArraySlice_l166_165 = (_zz_when_ArraySlice_l166_165 <= _zz_when_ArraySlice_l166_165_2);
  assign _zz_when_ArraySlice_l112_165 = (wReg % _zz__zz_when_ArraySlice_l112_165);
  assign when_ArraySlice_l112_165 = (_zz_when_ArraySlice_l112_165 != 6'h0);
  assign when_ArraySlice_l113_165 = (7'h40 <= _zz_when_ArraySlice_l113_165);
  always @(*) begin
    if(when_ArraySlice_l112_165) begin
      if(when_ArraySlice_l113_165) begin
        _zz_when_ArraySlice_l173_165 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_165 = (_zz__zz_when_ArraySlice_l173_165 - _zz__zz_when_ArraySlice_l173_165_3);
      end
    end else begin
      if(when_ArraySlice_l118_165) begin
        _zz_when_ArraySlice_l173_165 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_165 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_165 = (_zz_when_ArraySlice_l118_165 <= wReg);
  assign when_ArraySlice_l173_165 = (_zz_when_ArraySlice_l173_165_1 <= _zz_when_ArraySlice_l173_165_3);
  assign when_ArraySlice_l165_166 = (_zz_when_ArraySlice_l165_166 <= selectWriteFifo);
  assign when_ArraySlice_l166_166 = (_zz_when_ArraySlice_l166_166 <= _zz_when_ArraySlice_l166_166_2);
  assign _zz_when_ArraySlice_l112_166 = (wReg % _zz__zz_when_ArraySlice_l112_166);
  assign when_ArraySlice_l112_166 = (_zz_when_ArraySlice_l112_166 != 6'h0);
  assign when_ArraySlice_l113_166 = (7'h40 <= _zz_when_ArraySlice_l113_166);
  always @(*) begin
    if(when_ArraySlice_l112_166) begin
      if(when_ArraySlice_l113_166) begin
        _zz_when_ArraySlice_l173_166 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_166 = (_zz__zz_when_ArraySlice_l173_166 - _zz__zz_when_ArraySlice_l173_166_3);
      end
    end else begin
      if(when_ArraySlice_l118_166) begin
        _zz_when_ArraySlice_l173_166 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_166 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_166 = (_zz_when_ArraySlice_l118_166 <= wReg);
  assign when_ArraySlice_l173_166 = (_zz_when_ArraySlice_l173_166_1 <= _zz_when_ArraySlice_l173_166_3);
  assign when_ArraySlice_l165_167 = (_zz_when_ArraySlice_l165_167 <= selectWriteFifo);
  assign when_ArraySlice_l166_167 = (_zz_when_ArraySlice_l166_167 <= _zz_when_ArraySlice_l166_167_2);
  assign _zz_when_ArraySlice_l112_167 = (wReg % _zz__zz_when_ArraySlice_l112_167);
  assign when_ArraySlice_l112_167 = (_zz_when_ArraySlice_l112_167 != 6'h0);
  assign when_ArraySlice_l113_167 = (7'h40 <= _zz_when_ArraySlice_l113_167);
  always @(*) begin
    if(when_ArraySlice_l112_167) begin
      if(when_ArraySlice_l113_167) begin
        _zz_when_ArraySlice_l173_167 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_167 = (_zz__zz_when_ArraySlice_l173_167 - _zz__zz_when_ArraySlice_l173_167_3);
      end
    end else begin
      if(when_ArraySlice_l118_167) begin
        _zz_when_ArraySlice_l173_167 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_167 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_167 = (_zz_when_ArraySlice_l118_167 <= wReg);
  assign when_ArraySlice_l173_167 = (_zz_when_ArraySlice_l173_167_1 <= _zz_when_ArraySlice_l173_167_3);
  assign when_ArraySlice_l418_6 = (! ((((((_zz_when_ArraySlice_l418_6 && _zz_when_ArraySlice_l418_6_1) && (holdReadOp_4 == _zz_when_ArraySlice_l418_6_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l418_6_3 && _zz_when_ArraySlice_l418_6_4) && (debug_4_20 == _zz_when_ArraySlice_l418_6_5)) && (debug_5_20 == 1'b1)) && (debug_6_20 == 1'b1)) && (debug_7_20 == 1'b1))));
  assign when_ArraySlice_l421_6 = (wReg <= _zz_when_ArraySlice_l421_6_1);
  assign outputStreamArrayData_6_fire_3 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l425_6 = ((_zz_when_ArraySlice_l425_6 == 13'h0) && outputStreamArrayData_6_fire_3);
  assign outputStreamArrayData_6_fire_4 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l436_6 = ((handshakeTimes_6_value == _zz_when_ArraySlice_l436_6) && outputStreamArrayData_6_fire_4);
  assign _zz_when_ArraySlice_l94_20 = (hReg % _zz__zz_when_ArraySlice_l94_20);
  assign when_ArraySlice_l94_20 = (_zz_when_ArraySlice_l94_20 != 6'h0);
  assign when_ArraySlice_l95_20 = (7'h40 <= _zz_when_ArraySlice_l95_20);
  always @(*) begin
    if(when_ArraySlice_l94_20) begin
      if(when_ArraySlice_l95_20) begin
        _zz_when_ArraySlice_l437_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_6 = (_zz__zz_when_ArraySlice_l437_6 - _zz__zz_when_ArraySlice_l437_6_3);
      end
    end else begin
      if(when_ArraySlice_l99_20) begin
        _zz_when_ArraySlice_l437_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_6 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_20 = (_zz_when_ArraySlice_l99_20 <= hReg);
  assign when_ArraySlice_l437_6 = (_zz_when_ArraySlice_l437_6_1 < _zz_when_ArraySlice_l437_6_4);
  always @(*) begin
    debug_0_21 = 1'b0;
    if(when_ArraySlice_l165_168) begin
      if(when_ArraySlice_l166_168) begin
        debug_0_21 = 1'b1;
      end else begin
        debug_0_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_168) begin
        debug_0_21 = 1'b1;
      end else begin
        debug_0_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_21 = 1'b0;
    if(when_ArraySlice_l165_169) begin
      if(when_ArraySlice_l166_169) begin
        debug_1_21 = 1'b1;
      end else begin
        debug_1_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_169) begin
        debug_1_21 = 1'b1;
      end else begin
        debug_1_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_21 = 1'b0;
    if(when_ArraySlice_l165_170) begin
      if(when_ArraySlice_l166_170) begin
        debug_2_21 = 1'b1;
      end else begin
        debug_2_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_170) begin
        debug_2_21 = 1'b1;
      end else begin
        debug_2_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_21 = 1'b0;
    if(when_ArraySlice_l165_171) begin
      if(when_ArraySlice_l166_171) begin
        debug_3_21 = 1'b1;
      end else begin
        debug_3_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_171) begin
        debug_3_21 = 1'b1;
      end else begin
        debug_3_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_21 = 1'b0;
    if(when_ArraySlice_l165_172) begin
      if(when_ArraySlice_l166_172) begin
        debug_4_21 = 1'b1;
      end else begin
        debug_4_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_172) begin
        debug_4_21 = 1'b1;
      end else begin
        debug_4_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_21 = 1'b0;
    if(when_ArraySlice_l165_173) begin
      if(when_ArraySlice_l166_173) begin
        debug_5_21 = 1'b1;
      end else begin
        debug_5_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_173) begin
        debug_5_21 = 1'b1;
      end else begin
        debug_5_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_21 = 1'b0;
    if(when_ArraySlice_l165_174) begin
      if(when_ArraySlice_l166_174) begin
        debug_6_21 = 1'b1;
      end else begin
        debug_6_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_174) begin
        debug_6_21 = 1'b1;
      end else begin
        debug_6_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_21 = 1'b0;
    if(when_ArraySlice_l165_175) begin
      if(when_ArraySlice_l166_175) begin
        debug_7_21 = 1'b1;
      end else begin
        debug_7_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_175) begin
        debug_7_21 = 1'b1;
      end else begin
        debug_7_21 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_168 = (_zz_when_ArraySlice_l165_168 <= selectWriteFifo);
  assign when_ArraySlice_l166_168 = (_zz_when_ArraySlice_l166_168 <= _zz_when_ArraySlice_l166_168_1);
  assign _zz_when_ArraySlice_l112_168 = (wReg % _zz__zz_when_ArraySlice_l112_168);
  assign when_ArraySlice_l112_168 = (_zz_when_ArraySlice_l112_168 != 6'h0);
  assign when_ArraySlice_l113_168 = (7'h40 <= _zz_when_ArraySlice_l113_168);
  always @(*) begin
    if(when_ArraySlice_l112_168) begin
      if(when_ArraySlice_l113_168) begin
        _zz_when_ArraySlice_l173_168 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_168 = (_zz__zz_when_ArraySlice_l173_168 - _zz__zz_when_ArraySlice_l173_168_3);
      end
    end else begin
      if(when_ArraySlice_l118_168) begin
        _zz_when_ArraySlice_l173_168 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_168 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_168 = (_zz_when_ArraySlice_l118_168 <= wReg);
  assign when_ArraySlice_l173_168 = (_zz_when_ArraySlice_l173_168_1 <= _zz_when_ArraySlice_l173_168_2);
  assign when_ArraySlice_l165_169 = (_zz_when_ArraySlice_l165_169 <= selectWriteFifo);
  assign when_ArraySlice_l166_169 = (_zz_when_ArraySlice_l166_169 <= _zz_when_ArraySlice_l166_169_1);
  assign _zz_when_ArraySlice_l112_169 = (wReg % _zz__zz_when_ArraySlice_l112_169);
  assign when_ArraySlice_l112_169 = (_zz_when_ArraySlice_l112_169 != 6'h0);
  assign when_ArraySlice_l113_169 = (7'h40 <= _zz_when_ArraySlice_l113_169);
  always @(*) begin
    if(when_ArraySlice_l112_169) begin
      if(when_ArraySlice_l113_169) begin
        _zz_when_ArraySlice_l173_169 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_169 = (_zz__zz_when_ArraySlice_l173_169 - _zz__zz_when_ArraySlice_l173_169_3);
      end
    end else begin
      if(when_ArraySlice_l118_169) begin
        _zz_when_ArraySlice_l173_169 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_169 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_169 = (_zz_when_ArraySlice_l118_169 <= wReg);
  assign when_ArraySlice_l173_169 = (_zz_when_ArraySlice_l173_169_1 <= _zz_when_ArraySlice_l173_169_3);
  assign when_ArraySlice_l165_170 = (_zz_when_ArraySlice_l165_170 <= selectWriteFifo);
  assign when_ArraySlice_l166_170 = (_zz_when_ArraySlice_l166_170 <= _zz_when_ArraySlice_l166_170_1);
  assign _zz_when_ArraySlice_l112_170 = (wReg % _zz__zz_when_ArraySlice_l112_170);
  assign when_ArraySlice_l112_170 = (_zz_when_ArraySlice_l112_170 != 6'h0);
  assign when_ArraySlice_l113_170 = (7'h40 <= _zz_when_ArraySlice_l113_170);
  always @(*) begin
    if(when_ArraySlice_l112_170) begin
      if(when_ArraySlice_l113_170) begin
        _zz_when_ArraySlice_l173_170 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_170 = (_zz__zz_when_ArraySlice_l173_170 - _zz__zz_when_ArraySlice_l173_170_3);
      end
    end else begin
      if(when_ArraySlice_l118_170) begin
        _zz_when_ArraySlice_l173_170 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_170 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_170 = (_zz_when_ArraySlice_l118_170 <= wReg);
  assign when_ArraySlice_l173_170 = (_zz_when_ArraySlice_l173_170_1 <= _zz_when_ArraySlice_l173_170_3);
  assign when_ArraySlice_l165_171 = (_zz_when_ArraySlice_l165_171 <= selectWriteFifo);
  assign when_ArraySlice_l166_171 = (_zz_when_ArraySlice_l166_171 <= _zz_when_ArraySlice_l166_171_1);
  assign _zz_when_ArraySlice_l112_171 = (wReg % _zz__zz_when_ArraySlice_l112_171);
  assign when_ArraySlice_l112_171 = (_zz_when_ArraySlice_l112_171 != 6'h0);
  assign when_ArraySlice_l113_171 = (7'h40 <= _zz_when_ArraySlice_l113_171);
  always @(*) begin
    if(when_ArraySlice_l112_171) begin
      if(when_ArraySlice_l113_171) begin
        _zz_when_ArraySlice_l173_171 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_171 = (_zz__zz_when_ArraySlice_l173_171 - _zz__zz_when_ArraySlice_l173_171_3);
      end
    end else begin
      if(when_ArraySlice_l118_171) begin
        _zz_when_ArraySlice_l173_171 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_171 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_171 = (_zz_when_ArraySlice_l118_171 <= wReg);
  assign when_ArraySlice_l173_171 = (_zz_when_ArraySlice_l173_171_1 <= _zz_when_ArraySlice_l173_171_3);
  assign when_ArraySlice_l165_172 = (_zz_when_ArraySlice_l165_172 <= selectWriteFifo);
  assign when_ArraySlice_l166_172 = (_zz_when_ArraySlice_l166_172 <= _zz_when_ArraySlice_l166_172_1);
  assign _zz_when_ArraySlice_l112_172 = (wReg % _zz__zz_when_ArraySlice_l112_172);
  assign when_ArraySlice_l112_172 = (_zz_when_ArraySlice_l112_172 != 6'h0);
  assign when_ArraySlice_l113_172 = (7'h40 <= _zz_when_ArraySlice_l113_172);
  always @(*) begin
    if(when_ArraySlice_l112_172) begin
      if(when_ArraySlice_l113_172) begin
        _zz_when_ArraySlice_l173_172 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_172 = (_zz__zz_when_ArraySlice_l173_172 - _zz__zz_when_ArraySlice_l173_172_3);
      end
    end else begin
      if(when_ArraySlice_l118_172) begin
        _zz_when_ArraySlice_l173_172 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_172 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_172 = (_zz_when_ArraySlice_l118_172 <= wReg);
  assign when_ArraySlice_l173_172 = (_zz_when_ArraySlice_l173_172_1 <= _zz_when_ArraySlice_l173_172_3);
  assign when_ArraySlice_l165_173 = (_zz_when_ArraySlice_l165_173 <= selectWriteFifo);
  assign when_ArraySlice_l166_173 = (_zz_when_ArraySlice_l166_173 <= _zz_when_ArraySlice_l166_173_2);
  assign _zz_when_ArraySlice_l112_173 = (wReg % _zz__zz_when_ArraySlice_l112_173);
  assign when_ArraySlice_l112_173 = (_zz_when_ArraySlice_l112_173 != 6'h0);
  assign when_ArraySlice_l113_173 = (7'h40 <= _zz_when_ArraySlice_l113_173);
  always @(*) begin
    if(when_ArraySlice_l112_173) begin
      if(when_ArraySlice_l113_173) begin
        _zz_when_ArraySlice_l173_173 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_173 = (_zz__zz_when_ArraySlice_l173_173 - _zz__zz_when_ArraySlice_l173_173_3);
      end
    end else begin
      if(when_ArraySlice_l118_173) begin
        _zz_when_ArraySlice_l173_173 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_173 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_173 = (_zz_when_ArraySlice_l118_173 <= wReg);
  assign when_ArraySlice_l173_173 = (_zz_when_ArraySlice_l173_173_1 <= _zz_when_ArraySlice_l173_173_3);
  assign when_ArraySlice_l165_174 = (_zz_when_ArraySlice_l165_174 <= selectWriteFifo);
  assign when_ArraySlice_l166_174 = (_zz_when_ArraySlice_l166_174 <= _zz_when_ArraySlice_l166_174_2);
  assign _zz_when_ArraySlice_l112_174 = (wReg % _zz__zz_when_ArraySlice_l112_174);
  assign when_ArraySlice_l112_174 = (_zz_when_ArraySlice_l112_174 != 6'h0);
  assign when_ArraySlice_l113_174 = (7'h40 <= _zz_when_ArraySlice_l113_174);
  always @(*) begin
    if(when_ArraySlice_l112_174) begin
      if(when_ArraySlice_l113_174) begin
        _zz_when_ArraySlice_l173_174 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_174 = (_zz__zz_when_ArraySlice_l173_174 - _zz__zz_when_ArraySlice_l173_174_3);
      end
    end else begin
      if(when_ArraySlice_l118_174) begin
        _zz_when_ArraySlice_l173_174 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_174 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_174 = (_zz_when_ArraySlice_l118_174 <= wReg);
  assign when_ArraySlice_l173_174 = (_zz_when_ArraySlice_l173_174_1 <= _zz_when_ArraySlice_l173_174_3);
  assign when_ArraySlice_l165_175 = (_zz_when_ArraySlice_l165_175 <= selectWriteFifo);
  assign when_ArraySlice_l166_175 = (_zz_when_ArraySlice_l166_175 <= _zz_when_ArraySlice_l166_175_2);
  assign _zz_when_ArraySlice_l112_175 = (wReg % _zz__zz_when_ArraySlice_l112_175);
  assign when_ArraySlice_l112_175 = (_zz_when_ArraySlice_l112_175 != 6'h0);
  assign when_ArraySlice_l113_175 = (7'h40 <= _zz_when_ArraySlice_l113_175);
  always @(*) begin
    if(when_ArraySlice_l112_175) begin
      if(when_ArraySlice_l113_175) begin
        _zz_when_ArraySlice_l173_175 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_175 = (_zz__zz_when_ArraySlice_l173_175 - _zz__zz_when_ArraySlice_l173_175_3);
      end
    end else begin
      if(when_ArraySlice_l118_175) begin
        _zz_when_ArraySlice_l173_175 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_175 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_175 = (_zz_when_ArraySlice_l118_175 <= wReg);
  assign when_ArraySlice_l173_175 = (_zz_when_ArraySlice_l173_175_1 <= _zz_when_ArraySlice_l173_175_3);
  assign when_ArraySlice_l444_6 = (! ((((((_zz_when_ArraySlice_l444_6 && _zz_when_ArraySlice_l444_6_1) && (holdReadOp_4 == _zz_when_ArraySlice_l444_6_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l444_6_3 && _zz_when_ArraySlice_l444_6_4) && (debug_4_21 == _zz_when_ArraySlice_l444_6_5)) && (debug_5_21 == 1'b1)) && (debug_6_21 == 1'b1)) && (debug_7_21 == 1'b1))));
  assign outputStreamArrayData_6_fire_5 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l448_6 = ((_zz_when_ArraySlice_l448_6 == 13'h0) && outputStreamArrayData_6_fire_5);
  assign when_ArraySlice_l434_6 = (allowPadding_6 && (wReg <= _zz_when_ArraySlice_l434_6));
  assign outputStreamArrayData_6_fire_6 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l455_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l455_6);
  assign when_ArraySlice_l373_7 = (_zz_when_ArraySlice_l373_7 < wReg);
  assign when_ArraySlice_l374_7 = ((! holdReadOp_7) && (_zz_when_ArraySlice_l374_7 != 7'h0));
  assign _zz_outputStreamArrayData_7_valid = (selectReadFifo_7 + _zz__zz_outputStreamArrayData_7_valid);
  assign _zz_10 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_7_valid);
  assign _zz_io_pop_ready_7 = outputStreamArrayData_7_ready;
  assign when_ArraySlice_l379_7 = (! holdReadOp_7);
  assign outputStreamArrayData_7_fire = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l380_7 = ((_zz_when_ArraySlice_l380_7 < _zz_when_ArraySlice_l380_7_2) && outputStreamArrayData_7_fire);
  assign when_ArraySlice_l381_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l381_7);
  assign when_ArraySlice_l384_7 = (_zz_when_ArraySlice_l384_7 == 13'h0);
  assign outputStreamArrayData_7_fire_1 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l389_7 = ((_zz_when_ArraySlice_l389_7 == _zz_when_ArraySlice_l389_7_3) && outputStreamArrayData_7_fire_1);
  assign when_ArraySlice_l390_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l390_7);
  assign _zz_when_ArraySlice_l94_21 = (hReg % _zz__zz_when_ArraySlice_l94_21);
  assign when_ArraySlice_l94_21 = (_zz_when_ArraySlice_l94_21 != 6'h0);
  assign when_ArraySlice_l95_21 = (7'h40 <= _zz_when_ArraySlice_l95_21);
  always @(*) begin
    if(when_ArraySlice_l94_21) begin
      if(when_ArraySlice_l95_21) begin
        _zz_when_ArraySlice_l392_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_7 = (_zz__zz_when_ArraySlice_l392_7 - _zz__zz_when_ArraySlice_l392_7_3);
      end
    end else begin
      if(when_ArraySlice_l99_21) begin
        _zz_when_ArraySlice_l392_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l392_7 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_21 = (_zz_when_ArraySlice_l99_21 <= hReg);
  assign when_ArraySlice_l392_7 = (_zz_when_ArraySlice_l392_7_1 < _zz_when_ArraySlice_l392_7_4);
  always @(*) begin
    debug_0_22 = 1'b0;
    if(when_ArraySlice_l165_176) begin
      if(when_ArraySlice_l166_176) begin
        debug_0_22 = 1'b1;
      end else begin
        debug_0_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_176) begin
        debug_0_22 = 1'b1;
      end else begin
        debug_0_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_22 = 1'b0;
    if(when_ArraySlice_l165_177) begin
      if(when_ArraySlice_l166_177) begin
        debug_1_22 = 1'b1;
      end else begin
        debug_1_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_177) begin
        debug_1_22 = 1'b1;
      end else begin
        debug_1_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_22 = 1'b0;
    if(when_ArraySlice_l165_178) begin
      if(when_ArraySlice_l166_178) begin
        debug_2_22 = 1'b1;
      end else begin
        debug_2_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_178) begin
        debug_2_22 = 1'b1;
      end else begin
        debug_2_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_22 = 1'b0;
    if(when_ArraySlice_l165_179) begin
      if(when_ArraySlice_l166_179) begin
        debug_3_22 = 1'b1;
      end else begin
        debug_3_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_179) begin
        debug_3_22 = 1'b1;
      end else begin
        debug_3_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_22 = 1'b0;
    if(when_ArraySlice_l165_180) begin
      if(when_ArraySlice_l166_180) begin
        debug_4_22 = 1'b1;
      end else begin
        debug_4_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_180) begin
        debug_4_22 = 1'b1;
      end else begin
        debug_4_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_22 = 1'b0;
    if(when_ArraySlice_l165_181) begin
      if(when_ArraySlice_l166_181) begin
        debug_5_22 = 1'b1;
      end else begin
        debug_5_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_181) begin
        debug_5_22 = 1'b1;
      end else begin
        debug_5_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_22 = 1'b0;
    if(when_ArraySlice_l165_182) begin
      if(when_ArraySlice_l166_182) begin
        debug_6_22 = 1'b1;
      end else begin
        debug_6_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_182) begin
        debug_6_22 = 1'b1;
      end else begin
        debug_6_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_22 = 1'b0;
    if(when_ArraySlice_l165_183) begin
      if(when_ArraySlice_l166_183) begin
        debug_7_22 = 1'b1;
      end else begin
        debug_7_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_183) begin
        debug_7_22 = 1'b1;
      end else begin
        debug_7_22 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_176 = (_zz_when_ArraySlice_l165_176 <= selectWriteFifo);
  assign when_ArraySlice_l166_176 = (_zz_when_ArraySlice_l166_176 <= _zz_when_ArraySlice_l166_176_1);
  assign _zz_when_ArraySlice_l112_176 = (wReg % _zz__zz_when_ArraySlice_l112_176);
  assign when_ArraySlice_l112_176 = (_zz_when_ArraySlice_l112_176 != 6'h0);
  assign when_ArraySlice_l113_176 = (7'h40 <= _zz_when_ArraySlice_l113_176);
  always @(*) begin
    if(when_ArraySlice_l112_176) begin
      if(when_ArraySlice_l113_176) begin
        _zz_when_ArraySlice_l173_176 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_176 = (_zz__zz_when_ArraySlice_l173_176 - _zz__zz_when_ArraySlice_l173_176_3);
      end
    end else begin
      if(when_ArraySlice_l118_176) begin
        _zz_when_ArraySlice_l173_176 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_176 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_176 = (_zz_when_ArraySlice_l118_176 <= wReg);
  assign when_ArraySlice_l173_176 = (_zz_when_ArraySlice_l173_176_1 <= _zz_when_ArraySlice_l173_176_2);
  assign when_ArraySlice_l165_177 = (_zz_when_ArraySlice_l165_177 <= selectWriteFifo);
  assign when_ArraySlice_l166_177 = (_zz_when_ArraySlice_l166_177 <= _zz_when_ArraySlice_l166_177_1);
  assign _zz_when_ArraySlice_l112_177 = (wReg % _zz__zz_when_ArraySlice_l112_177);
  assign when_ArraySlice_l112_177 = (_zz_when_ArraySlice_l112_177 != 6'h0);
  assign when_ArraySlice_l113_177 = (7'h40 <= _zz_when_ArraySlice_l113_177);
  always @(*) begin
    if(when_ArraySlice_l112_177) begin
      if(when_ArraySlice_l113_177) begin
        _zz_when_ArraySlice_l173_177 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_177 = (_zz__zz_when_ArraySlice_l173_177 - _zz__zz_when_ArraySlice_l173_177_3);
      end
    end else begin
      if(when_ArraySlice_l118_177) begin
        _zz_when_ArraySlice_l173_177 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_177 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_177 = (_zz_when_ArraySlice_l118_177 <= wReg);
  assign when_ArraySlice_l173_177 = (_zz_when_ArraySlice_l173_177_1 <= _zz_when_ArraySlice_l173_177_3);
  assign when_ArraySlice_l165_178 = (_zz_when_ArraySlice_l165_178 <= selectWriteFifo);
  assign when_ArraySlice_l166_178 = (_zz_when_ArraySlice_l166_178 <= _zz_when_ArraySlice_l166_178_1);
  assign _zz_when_ArraySlice_l112_178 = (wReg % _zz__zz_when_ArraySlice_l112_178);
  assign when_ArraySlice_l112_178 = (_zz_when_ArraySlice_l112_178 != 6'h0);
  assign when_ArraySlice_l113_178 = (7'h40 <= _zz_when_ArraySlice_l113_178);
  always @(*) begin
    if(when_ArraySlice_l112_178) begin
      if(when_ArraySlice_l113_178) begin
        _zz_when_ArraySlice_l173_178 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_178 = (_zz__zz_when_ArraySlice_l173_178 - _zz__zz_when_ArraySlice_l173_178_3);
      end
    end else begin
      if(when_ArraySlice_l118_178) begin
        _zz_when_ArraySlice_l173_178 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_178 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_178 = (_zz_when_ArraySlice_l118_178 <= wReg);
  assign when_ArraySlice_l173_178 = (_zz_when_ArraySlice_l173_178_1 <= _zz_when_ArraySlice_l173_178_3);
  assign when_ArraySlice_l165_179 = (_zz_when_ArraySlice_l165_179 <= selectWriteFifo);
  assign when_ArraySlice_l166_179 = (_zz_when_ArraySlice_l166_179 <= _zz_when_ArraySlice_l166_179_1);
  assign _zz_when_ArraySlice_l112_179 = (wReg % _zz__zz_when_ArraySlice_l112_179);
  assign when_ArraySlice_l112_179 = (_zz_when_ArraySlice_l112_179 != 6'h0);
  assign when_ArraySlice_l113_179 = (7'h40 <= _zz_when_ArraySlice_l113_179);
  always @(*) begin
    if(when_ArraySlice_l112_179) begin
      if(when_ArraySlice_l113_179) begin
        _zz_when_ArraySlice_l173_179 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_179 = (_zz__zz_when_ArraySlice_l173_179 - _zz__zz_when_ArraySlice_l173_179_3);
      end
    end else begin
      if(when_ArraySlice_l118_179) begin
        _zz_when_ArraySlice_l173_179 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_179 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_179 = (_zz_when_ArraySlice_l118_179 <= wReg);
  assign when_ArraySlice_l173_179 = (_zz_when_ArraySlice_l173_179_1 <= _zz_when_ArraySlice_l173_179_3);
  assign when_ArraySlice_l165_180 = (_zz_when_ArraySlice_l165_180 <= selectWriteFifo);
  assign when_ArraySlice_l166_180 = (_zz_when_ArraySlice_l166_180 <= _zz_when_ArraySlice_l166_180_1);
  assign _zz_when_ArraySlice_l112_180 = (wReg % _zz__zz_when_ArraySlice_l112_180);
  assign when_ArraySlice_l112_180 = (_zz_when_ArraySlice_l112_180 != 6'h0);
  assign when_ArraySlice_l113_180 = (7'h40 <= _zz_when_ArraySlice_l113_180);
  always @(*) begin
    if(when_ArraySlice_l112_180) begin
      if(when_ArraySlice_l113_180) begin
        _zz_when_ArraySlice_l173_180 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_180 = (_zz__zz_when_ArraySlice_l173_180 - _zz__zz_when_ArraySlice_l173_180_3);
      end
    end else begin
      if(when_ArraySlice_l118_180) begin
        _zz_when_ArraySlice_l173_180 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_180 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_180 = (_zz_when_ArraySlice_l118_180 <= wReg);
  assign when_ArraySlice_l173_180 = (_zz_when_ArraySlice_l173_180_1 <= _zz_when_ArraySlice_l173_180_3);
  assign when_ArraySlice_l165_181 = (_zz_when_ArraySlice_l165_181 <= selectWriteFifo);
  assign when_ArraySlice_l166_181 = (_zz_when_ArraySlice_l166_181 <= _zz_when_ArraySlice_l166_181_2);
  assign _zz_when_ArraySlice_l112_181 = (wReg % _zz__zz_when_ArraySlice_l112_181);
  assign when_ArraySlice_l112_181 = (_zz_when_ArraySlice_l112_181 != 6'h0);
  assign when_ArraySlice_l113_181 = (7'h40 <= _zz_when_ArraySlice_l113_181);
  always @(*) begin
    if(when_ArraySlice_l112_181) begin
      if(when_ArraySlice_l113_181) begin
        _zz_when_ArraySlice_l173_181 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_181 = (_zz__zz_when_ArraySlice_l173_181 - _zz__zz_when_ArraySlice_l173_181_3);
      end
    end else begin
      if(when_ArraySlice_l118_181) begin
        _zz_when_ArraySlice_l173_181 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_181 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_181 = (_zz_when_ArraySlice_l118_181 <= wReg);
  assign when_ArraySlice_l173_181 = (_zz_when_ArraySlice_l173_181_1 <= _zz_when_ArraySlice_l173_181_3);
  assign when_ArraySlice_l165_182 = (_zz_when_ArraySlice_l165_182 <= selectWriteFifo);
  assign when_ArraySlice_l166_182 = (_zz_when_ArraySlice_l166_182 <= _zz_when_ArraySlice_l166_182_2);
  assign _zz_when_ArraySlice_l112_182 = (wReg % _zz__zz_when_ArraySlice_l112_182);
  assign when_ArraySlice_l112_182 = (_zz_when_ArraySlice_l112_182 != 6'h0);
  assign when_ArraySlice_l113_182 = (7'h40 <= _zz_when_ArraySlice_l113_182);
  always @(*) begin
    if(when_ArraySlice_l112_182) begin
      if(when_ArraySlice_l113_182) begin
        _zz_when_ArraySlice_l173_182 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_182 = (_zz__zz_when_ArraySlice_l173_182 - _zz__zz_when_ArraySlice_l173_182_3);
      end
    end else begin
      if(when_ArraySlice_l118_182) begin
        _zz_when_ArraySlice_l173_182 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_182 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_182 = (_zz_when_ArraySlice_l118_182 <= wReg);
  assign when_ArraySlice_l173_182 = (_zz_when_ArraySlice_l173_182_1 <= _zz_when_ArraySlice_l173_182_3);
  assign when_ArraySlice_l165_183 = (_zz_when_ArraySlice_l165_183 <= selectWriteFifo);
  assign when_ArraySlice_l166_183 = (_zz_when_ArraySlice_l166_183 <= _zz_when_ArraySlice_l166_183_2);
  assign _zz_when_ArraySlice_l112_183 = (wReg % _zz__zz_when_ArraySlice_l112_183);
  assign when_ArraySlice_l112_183 = (_zz_when_ArraySlice_l112_183 != 6'h0);
  assign when_ArraySlice_l113_183 = (7'h40 <= _zz_when_ArraySlice_l113_183);
  always @(*) begin
    if(when_ArraySlice_l112_183) begin
      if(when_ArraySlice_l113_183) begin
        _zz_when_ArraySlice_l173_183 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_183 = (_zz__zz_when_ArraySlice_l173_183 - _zz__zz_when_ArraySlice_l173_183_3);
      end
    end else begin
      if(when_ArraySlice_l118_183) begin
        _zz_when_ArraySlice_l173_183 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_183 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_183 = (_zz_when_ArraySlice_l118_183 <= wReg);
  assign when_ArraySlice_l173_183 = (_zz_when_ArraySlice_l173_183_1 <= _zz_when_ArraySlice_l173_183_3);
  assign when_ArraySlice_l398_7 = (! ((((((_zz_when_ArraySlice_l398_7_1 && _zz_when_ArraySlice_l398_7_2) && (holdReadOp_4 == _zz_when_ArraySlice_l398_7_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l398_7_4 && _zz_when_ArraySlice_l398_7_5) && (debug_4_22 == _zz_when_ArraySlice_l398_7_6)) && (debug_5_22 == 1'b1)) && (debug_6_22 == 1'b1)) && (debug_7_22 == 1'b1))));
  assign when_ArraySlice_l401_7 = (wReg <= _zz_when_ArraySlice_l401_7_1);
  assign when_ArraySlice_l405_7 = (_zz_when_ArraySlice_l405_7 == 13'h0);
  assign when_ArraySlice_l409_7 = (_zz_when_ArraySlice_l409_7 == 7'h0);
  assign outputStreamArrayData_7_fire_2 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l410_7 = ((handshakeTimes_7_value == _zz_when_ArraySlice_l410_7) && outputStreamArrayData_7_fire_2);
  assign _zz_when_ArraySlice_l94_22 = (hReg % _zz__zz_when_ArraySlice_l94_22);
  assign when_ArraySlice_l94_22 = (_zz_when_ArraySlice_l94_22 != 6'h0);
  assign when_ArraySlice_l95_22 = (7'h40 <= _zz_when_ArraySlice_l95_22);
  always @(*) begin
    if(when_ArraySlice_l94_22) begin
      if(when_ArraySlice_l95_22) begin
        _zz_when_ArraySlice_l412_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_7 = (_zz__zz_when_ArraySlice_l412_7 - _zz__zz_when_ArraySlice_l412_7_3);
      end
    end else begin
      if(when_ArraySlice_l99_22) begin
        _zz_when_ArraySlice_l412_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l412_7 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_22 = (_zz_when_ArraySlice_l99_22 <= hReg);
  assign when_ArraySlice_l412_7 = (_zz_when_ArraySlice_l412_7_1 < _zz_when_ArraySlice_l412_7_4);
  always @(*) begin
    debug_0_23 = 1'b0;
    if(when_ArraySlice_l165_184) begin
      if(when_ArraySlice_l166_184) begin
        debug_0_23 = 1'b1;
      end else begin
        debug_0_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_184) begin
        debug_0_23 = 1'b1;
      end else begin
        debug_0_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_23 = 1'b0;
    if(when_ArraySlice_l165_185) begin
      if(when_ArraySlice_l166_185) begin
        debug_1_23 = 1'b1;
      end else begin
        debug_1_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_185) begin
        debug_1_23 = 1'b1;
      end else begin
        debug_1_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_23 = 1'b0;
    if(when_ArraySlice_l165_186) begin
      if(when_ArraySlice_l166_186) begin
        debug_2_23 = 1'b1;
      end else begin
        debug_2_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_186) begin
        debug_2_23 = 1'b1;
      end else begin
        debug_2_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_23 = 1'b0;
    if(when_ArraySlice_l165_187) begin
      if(when_ArraySlice_l166_187) begin
        debug_3_23 = 1'b1;
      end else begin
        debug_3_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_187) begin
        debug_3_23 = 1'b1;
      end else begin
        debug_3_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_23 = 1'b0;
    if(when_ArraySlice_l165_188) begin
      if(when_ArraySlice_l166_188) begin
        debug_4_23 = 1'b1;
      end else begin
        debug_4_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_188) begin
        debug_4_23 = 1'b1;
      end else begin
        debug_4_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_23 = 1'b0;
    if(when_ArraySlice_l165_189) begin
      if(when_ArraySlice_l166_189) begin
        debug_5_23 = 1'b1;
      end else begin
        debug_5_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_189) begin
        debug_5_23 = 1'b1;
      end else begin
        debug_5_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_23 = 1'b0;
    if(when_ArraySlice_l165_190) begin
      if(when_ArraySlice_l166_190) begin
        debug_6_23 = 1'b1;
      end else begin
        debug_6_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_190) begin
        debug_6_23 = 1'b1;
      end else begin
        debug_6_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_23 = 1'b0;
    if(when_ArraySlice_l165_191) begin
      if(when_ArraySlice_l166_191) begin
        debug_7_23 = 1'b1;
      end else begin
        debug_7_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_191) begin
        debug_7_23 = 1'b1;
      end else begin
        debug_7_23 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_184 = (_zz_when_ArraySlice_l165_184 <= selectWriteFifo);
  assign when_ArraySlice_l166_184 = (_zz_when_ArraySlice_l166_184 <= _zz_when_ArraySlice_l166_184_1);
  assign _zz_when_ArraySlice_l112_184 = (wReg % _zz__zz_when_ArraySlice_l112_184);
  assign when_ArraySlice_l112_184 = (_zz_when_ArraySlice_l112_184 != 6'h0);
  assign when_ArraySlice_l113_184 = (7'h40 <= _zz_when_ArraySlice_l113_184);
  always @(*) begin
    if(when_ArraySlice_l112_184) begin
      if(when_ArraySlice_l113_184) begin
        _zz_when_ArraySlice_l173_184 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_184 = (_zz__zz_when_ArraySlice_l173_184 - _zz__zz_when_ArraySlice_l173_184_3);
      end
    end else begin
      if(when_ArraySlice_l118_184) begin
        _zz_when_ArraySlice_l173_184 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_184 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_184 = (_zz_when_ArraySlice_l118_184 <= wReg);
  assign when_ArraySlice_l173_184 = (_zz_when_ArraySlice_l173_184_1 <= _zz_when_ArraySlice_l173_184_2);
  assign when_ArraySlice_l165_185 = (_zz_when_ArraySlice_l165_185 <= selectWriteFifo);
  assign when_ArraySlice_l166_185 = (_zz_when_ArraySlice_l166_185 <= _zz_when_ArraySlice_l166_185_1);
  assign _zz_when_ArraySlice_l112_185 = (wReg % _zz__zz_when_ArraySlice_l112_185);
  assign when_ArraySlice_l112_185 = (_zz_when_ArraySlice_l112_185 != 6'h0);
  assign when_ArraySlice_l113_185 = (7'h40 <= _zz_when_ArraySlice_l113_185);
  always @(*) begin
    if(when_ArraySlice_l112_185) begin
      if(when_ArraySlice_l113_185) begin
        _zz_when_ArraySlice_l173_185 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_185 = (_zz__zz_when_ArraySlice_l173_185 - _zz__zz_when_ArraySlice_l173_185_3);
      end
    end else begin
      if(when_ArraySlice_l118_185) begin
        _zz_when_ArraySlice_l173_185 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_185 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_185 = (_zz_when_ArraySlice_l118_185 <= wReg);
  assign when_ArraySlice_l173_185 = (_zz_when_ArraySlice_l173_185_1 <= _zz_when_ArraySlice_l173_185_3);
  assign when_ArraySlice_l165_186 = (_zz_when_ArraySlice_l165_186 <= selectWriteFifo);
  assign when_ArraySlice_l166_186 = (_zz_when_ArraySlice_l166_186 <= _zz_when_ArraySlice_l166_186_1);
  assign _zz_when_ArraySlice_l112_186 = (wReg % _zz__zz_when_ArraySlice_l112_186);
  assign when_ArraySlice_l112_186 = (_zz_when_ArraySlice_l112_186 != 6'h0);
  assign when_ArraySlice_l113_186 = (7'h40 <= _zz_when_ArraySlice_l113_186);
  always @(*) begin
    if(when_ArraySlice_l112_186) begin
      if(when_ArraySlice_l113_186) begin
        _zz_when_ArraySlice_l173_186 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_186 = (_zz__zz_when_ArraySlice_l173_186 - _zz__zz_when_ArraySlice_l173_186_3);
      end
    end else begin
      if(when_ArraySlice_l118_186) begin
        _zz_when_ArraySlice_l173_186 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_186 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_186 = (_zz_when_ArraySlice_l118_186 <= wReg);
  assign when_ArraySlice_l173_186 = (_zz_when_ArraySlice_l173_186_1 <= _zz_when_ArraySlice_l173_186_3);
  assign when_ArraySlice_l165_187 = (_zz_when_ArraySlice_l165_187 <= selectWriteFifo);
  assign when_ArraySlice_l166_187 = (_zz_when_ArraySlice_l166_187 <= _zz_when_ArraySlice_l166_187_1);
  assign _zz_when_ArraySlice_l112_187 = (wReg % _zz__zz_when_ArraySlice_l112_187);
  assign when_ArraySlice_l112_187 = (_zz_when_ArraySlice_l112_187 != 6'h0);
  assign when_ArraySlice_l113_187 = (7'h40 <= _zz_when_ArraySlice_l113_187);
  always @(*) begin
    if(when_ArraySlice_l112_187) begin
      if(when_ArraySlice_l113_187) begin
        _zz_when_ArraySlice_l173_187 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_187 = (_zz__zz_when_ArraySlice_l173_187 - _zz__zz_when_ArraySlice_l173_187_3);
      end
    end else begin
      if(when_ArraySlice_l118_187) begin
        _zz_when_ArraySlice_l173_187 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_187 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_187 = (_zz_when_ArraySlice_l118_187 <= wReg);
  assign when_ArraySlice_l173_187 = (_zz_when_ArraySlice_l173_187_1 <= _zz_when_ArraySlice_l173_187_3);
  assign when_ArraySlice_l165_188 = (_zz_when_ArraySlice_l165_188 <= selectWriteFifo);
  assign when_ArraySlice_l166_188 = (_zz_when_ArraySlice_l166_188 <= _zz_when_ArraySlice_l166_188_1);
  assign _zz_when_ArraySlice_l112_188 = (wReg % _zz__zz_when_ArraySlice_l112_188);
  assign when_ArraySlice_l112_188 = (_zz_when_ArraySlice_l112_188 != 6'h0);
  assign when_ArraySlice_l113_188 = (7'h40 <= _zz_when_ArraySlice_l113_188);
  always @(*) begin
    if(when_ArraySlice_l112_188) begin
      if(when_ArraySlice_l113_188) begin
        _zz_when_ArraySlice_l173_188 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_188 = (_zz__zz_when_ArraySlice_l173_188 - _zz__zz_when_ArraySlice_l173_188_3);
      end
    end else begin
      if(when_ArraySlice_l118_188) begin
        _zz_when_ArraySlice_l173_188 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_188 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_188 = (_zz_when_ArraySlice_l118_188 <= wReg);
  assign when_ArraySlice_l173_188 = (_zz_when_ArraySlice_l173_188_1 <= _zz_when_ArraySlice_l173_188_3);
  assign when_ArraySlice_l165_189 = (_zz_when_ArraySlice_l165_189 <= selectWriteFifo);
  assign when_ArraySlice_l166_189 = (_zz_when_ArraySlice_l166_189 <= _zz_when_ArraySlice_l166_189_2);
  assign _zz_when_ArraySlice_l112_189 = (wReg % _zz__zz_when_ArraySlice_l112_189);
  assign when_ArraySlice_l112_189 = (_zz_when_ArraySlice_l112_189 != 6'h0);
  assign when_ArraySlice_l113_189 = (7'h40 <= _zz_when_ArraySlice_l113_189);
  always @(*) begin
    if(when_ArraySlice_l112_189) begin
      if(when_ArraySlice_l113_189) begin
        _zz_when_ArraySlice_l173_189 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_189 = (_zz__zz_when_ArraySlice_l173_189 - _zz__zz_when_ArraySlice_l173_189_3);
      end
    end else begin
      if(when_ArraySlice_l118_189) begin
        _zz_when_ArraySlice_l173_189 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_189 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_189 = (_zz_when_ArraySlice_l118_189 <= wReg);
  assign when_ArraySlice_l173_189 = (_zz_when_ArraySlice_l173_189_1 <= _zz_when_ArraySlice_l173_189_3);
  assign when_ArraySlice_l165_190 = (_zz_when_ArraySlice_l165_190 <= selectWriteFifo);
  assign when_ArraySlice_l166_190 = (_zz_when_ArraySlice_l166_190 <= _zz_when_ArraySlice_l166_190_2);
  assign _zz_when_ArraySlice_l112_190 = (wReg % _zz__zz_when_ArraySlice_l112_190);
  assign when_ArraySlice_l112_190 = (_zz_when_ArraySlice_l112_190 != 6'h0);
  assign when_ArraySlice_l113_190 = (7'h40 <= _zz_when_ArraySlice_l113_190);
  always @(*) begin
    if(when_ArraySlice_l112_190) begin
      if(when_ArraySlice_l113_190) begin
        _zz_when_ArraySlice_l173_190 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_190 = (_zz__zz_when_ArraySlice_l173_190 - _zz__zz_when_ArraySlice_l173_190_3);
      end
    end else begin
      if(when_ArraySlice_l118_190) begin
        _zz_when_ArraySlice_l173_190 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_190 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_190 = (_zz_when_ArraySlice_l118_190 <= wReg);
  assign when_ArraySlice_l173_190 = (_zz_when_ArraySlice_l173_190_1 <= _zz_when_ArraySlice_l173_190_3);
  assign when_ArraySlice_l165_191 = (_zz_when_ArraySlice_l165_191 <= selectWriteFifo);
  assign when_ArraySlice_l166_191 = (_zz_when_ArraySlice_l166_191 <= _zz_when_ArraySlice_l166_191_2);
  assign _zz_when_ArraySlice_l112_191 = (wReg % _zz__zz_when_ArraySlice_l112_191);
  assign when_ArraySlice_l112_191 = (_zz_when_ArraySlice_l112_191 != 6'h0);
  assign when_ArraySlice_l113_191 = (7'h40 <= _zz_when_ArraySlice_l113_191);
  always @(*) begin
    if(when_ArraySlice_l112_191) begin
      if(when_ArraySlice_l113_191) begin
        _zz_when_ArraySlice_l173_191 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_191 = (_zz__zz_when_ArraySlice_l173_191 - _zz__zz_when_ArraySlice_l173_191_3);
      end
    end else begin
      if(when_ArraySlice_l118_191) begin
        _zz_when_ArraySlice_l173_191 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_191 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_191 = (_zz_when_ArraySlice_l118_191 <= wReg);
  assign when_ArraySlice_l173_191 = (_zz_when_ArraySlice_l173_191_1 <= _zz_when_ArraySlice_l173_191_3);
  assign when_ArraySlice_l418_7 = (! ((((((_zz_when_ArraySlice_l418_7 && _zz_when_ArraySlice_l418_7_1) && (holdReadOp_4 == _zz_when_ArraySlice_l418_7_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l418_7_3 && _zz_when_ArraySlice_l418_7_4) && (debug_4_23 == _zz_when_ArraySlice_l418_7_5)) && (debug_5_23 == 1'b1)) && (debug_6_23 == 1'b1)) && (debug_7_23 == 1'b1))));
  assign when_ArraySlice_l421_7 = (wReg <= _zz_when_ArraySlice_l421_7_1);
  assign outputStreamArrayData_7_fire_3 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l425_7 = ((_zz_when_ArraySlice_l425_7 == 13'h0) && outputStreamArrayData_7_fire_3);
  assign outputStreamArrayData_7_fire_4 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l436_7 = ((handshakeTimes_7_value == _zz_when_ArraySlice_l436_7) && outputStreamArrayData_7_fire_4);
  assign _zz_when_ArraySlice_l94_23 = (hReg % _zz__zz_when_ArraySlice_l94_23);
  assign when_ArraySlice_l94_23 = (_zz_when_ArraySlice_l94_23 != 6'h0);
  assign when_ArraySlice_l95_23 = (7'h40 <= _zz_when_ArraySlice_l95_23);
  always @(*) begin
    if(when_ArraySlice_l94_23) begin
      if(when_ArraySlice_l95_23) begin
        _zz_when_ArraySlice_l437_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_7 = (_zz__zz_when_ArraySlice_l437_7 - _zz__zz_when_ArraySlice_l437_7_3);
      end
    end else begin
      if(when_ArraySlice_l99_23) begin
        _zz_when_ArraySlice_l437_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l437_7 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_23 = (_zz_when_ArraySlice_l99_23 <= hReg);
  assign when_ArraySlice_l437_7 = (_zz_when_ArraySlice_l437_7_1 < _zz_when_ArraySlice_l437_7_4);
  always @(*) begin
    debug_0_24 = 1'b0;
    if(when_ArraySlice_l165_192) begin
      if(when_ArraySlice_l166_192) begin
        debug_0_24 = 1'b1;
      end else begin
        debug_0_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_192) begin
        debug_0_24 = 1'b1;
      end else begin
        debug_0_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_24 = 1'b0;
    if(when_ArraySlice_l165_193) begin
      if(when_ArraySlice_l166_193) begin
        debug_1_24 = 1'b1;
      end else begin
        debug_1_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_193) begin
        debug_1_24 = 1'b1;
      end else begin
        debug_1_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_24 = 1'b0;
    if(when_ArraySlice_l165_194) begin
      if(when_ArraySlice_l166_194) begin
        debug_2_24 = 1'b1;
      end else begin
        debug_2_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_194) begin
        debug_2_24 = 1'b1;
      end else begin
        debug_2_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_24 = 1'b0;
    if(when_ArraySlice_l165_195) begin
      if(when_ArraySlice_l166_195) begin
        debug_3_24 = 1'b1;
      end else begin
        debug_3_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_195) begin
        debug_3_24 = 1'b1;
      end else begin
        debug_3_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_24 = 1'b0;
    if(when_ArraySlice_l165_196) begin
      if(when_ArraySlice_l166_196) begin
        debug_4_24 = 1'b1;
      end else begin
        debug_4_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_196) begin
        debug_4_24 = 1'b1;
      end else begin
        debug_4_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_24 = 1'b0;
    if(when_ArraySlice_l165_197) begin
      if(when_ArraySlice_l166_197) begin
        debug_5_24 = 1'b1;
      end else begin
        debug_5_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_197) begin
        debug_5_24 = 1'b1;
      end else begin
        debug_5_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_24 = 1'b0;
    if(when_ArraySlice_l165_198) begin
      if(when_ArraySlice_l166_198) begin
        debug_6_24 = 1'b1;
      end else begin
        debug_6_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_198) begin
        debug_6_24 = 1'b1;
      end else begin
        debug_6_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_24 = 1'b0;
    if(when_ArraySlice_l165_199) begin
      if(when_ArraySlice_l166_199) begin
        debug_7_24 = 1'b1;
      end else begin
        debug_7_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_199) begin
        debug_7_24 = 1'b1;
      end else begin
        debug_7_24 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_192 = (_zz_when_ArraySlice_l165_192 <= selectWriteFifo);
  assign when_ArraySlice_l166_192 = (_zz_when_ArraySlice_l166_192 <= _zz_when_ArraySlice_l166_192_1);
  assign _zz_when_ArraySlice_l112_192 = (wReg % _zz__zz_when_ArraySlice_l112_192);
  assign when_ArraySlice_l112_192 = (_zz_when_ArraySlice_l112_192 != 6'h0);
  assign when_ArraySlice_l113_192 = (7'h40 <= _zz_when_ArraySlice_l113_192);
  always @(*) begin
    if(when_ArraySlice_l112_192) begin
      if(when_ArraySlice_l113_192) begin
        _zz_when_ArraySlice_l173_192 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_192 = (_zz__zz_when_ArraySlice_l173_192 - _zz__zz_when_ArraySlice_l173_192_3);
      end
    end else begin
      if(when_ArraySlice_l118_192) begin
        _zz_when_ArraySlice_l173_192 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_192 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_192 = (_zz_when_ArraySlice_l118_192 <= wReg);
  assign when_ArraySlice_l173_192 = (_zz_when_ArraySlice_l173_192_1 <= _zz_when_ArraySlice_l173_192_2);
  assign when_ArraySlice_l165_193 = (_zz_when_ArraySlice_l165_193 <= selectWriteFifo);
  assign when_ArraySlice_l166_193 = (_zz_when_ArraySlice_l166_193 <= _zz_when_ArraySlice_l166_193_1);
  assign _zz_when_ArraySlice_l112_193 = (wReg % _zz__zz_when_ArraySlice_l112_193);
  assign when_ArraySlice_l112_193 = (_zz_when_ArraySlice_l112_193 != 6'h0);
  assign when_ArraySlice_l113_193 = (7'h40 <= _zz_when_ArraySlice_l113_193);
  always @(*) begin
    if(when_ArraySlice_l112_193) begin
      if(when_ArraySlice_l113_193) begin
        _zz_when_ArraySlice_l173_193 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_193 = (_zz__zz_when_ArraySlice_l173_193 - _zz__zz_when_ArraySlice_l173_193_3);
      end
    end else begin
      if(when_ArraySlice_l118_193) begin
        _zz_when_ArraySlice_l173_193 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_193 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_193 = (_zz_when_ArraySlice_l118_193 <= wReg);
  assign when_ArraySlice_l173_193 = (_zz_when_ArraySlice_l173_193_1 <= _zz_when_ArraySlice_l173_193_3);
  assign when_ArraySlice_l165_194 = (_zz_when_ArraySlice_l165_194 <= selectWriteFifo);
  assign when_ArraySlice_l166_194 = (_zz_when_ArraySlice_l166_194 <= _zz_when_ArraySlice_l166_194_1);
  assign _zz_when_ArraySlice_l112_194 = (wReg % _zz__zz_when_ArraySlice_l112_194);
  assign when_ArraySlice_l112_194 = (_zz_when_ArraySlice_l112_194 != 6'h0);
  assign when_ArraySlice_l113_194 = (7'h40 <= _zz_when_ArraySlice_l113_194);
  always @(*) begin
    if(when_ArraySlice_l112_194) begin
      if(when_ArraySlice_l113_194) begin
        _zz_when_ArraySlice_l173_194 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_194 = (_zz__zz_when_ArraySlice_l173_194 - _zz__zz_when_ArraySlice_l173_194_3);
      end
    end else begin
      if(when_ArraySlice_l118_194) begin
        _zz_when_ArraySlice_l173_194 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_194 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_194 = (_zz_when_ArraySlice_l118_194 <= wReg);
  assign when_ArraySlice_l173_194 = (_zz_when_ArraySlice_l173_194_1 <= _zz_when_ArraySlice_l173_194_3);
  assign when_ArraySlice_l165_195 = (_zz_when_ArraySlice_l165_195 <= selectWriteFifo);
  assign when_ArraySlice_l166_195 = (_zz_when_ArraySlice_l166_195 <= _zz_when_ArraySlice_l166_195_1);
  assign _zz_when_ArraySlice_l112_195 = (wReg % _zz__zz_when_ArraySlice_l112_195);
  assign when_ArraySlice_l112_195 = (_zz_when_ArraySlice_l112_195 != 6'h0);
  assign when_ArraySlice_l113_195 = (7'h40 <= _zz_when_ArraySlice_l113_195);
  always @(*) begin
    if(when_ArraySlice_l112_195) begin
      if(when_ArraySlice_l113_195) begin
        _zz_when_ArraySlice_l173_195 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_195 = (_zz__zz_when_ArraySlice_l173_195 - _zz__zz_when_ArraySlice_l173_195_3);
      end
    end else begin
      if(when_ArraySlice_l118_195) begin
        _zz_when_ArraySlice_l173_195 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_195 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_195 = (_zz_when_ArraySlice_l118_195 <= wReg);
  assign when_ArraySlice_l173_195 = (_zz_when_ArraySlice_l173_195_1 <= _zz_when_ArraySlice_l173_195_3);
  assign when_ArraySlice_l165_196 = (_zz_when_ArraySlice_l165_196 <= selectWriteFifo);
  assign when_ArraySlice_l166_196 = (_zz_when_ArraySlice_l166_196 <= _zz_when_ArraySlice_l166_196_1);
  assign _zz_when_ArraySlice_l112_196 = (wReg % _zz__zz_when_ArraySlice_l112_196);
  assign when_ArraySlice_l112_196 = (_zz_when_ArraySlice_l112_196 != 6'h0);
  assign when_ArraySlice_l113_196 = (7'h40 <= _zz_when_ArraySlice_l113_196);
  always @(*) begin
    if(when_ArraySlice_l112_196) begin
      if(when_ArraySlice_l113_196) begin
        _zz_when_ArraySlice_l173_196 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_196 = (_zz__zz_when_ArraySlice_l173_196 - _zz__zz_when_ArraySlice_l173_196_3);
      end
    end else begin
      if(when_ArraySlice_l118_196) begin
        _zz_when_ArraySlice_l173_196 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_196 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_196 = (_zz_when_ArraySlice_l118_196 <= wReg);
  assign when_ArraySlice_l173_196 = (_zz_when_ArraySlice_l173_196_1 <= _zz_when_ArraySlice_l173_196_3);
  assign when_ArraySlice_l165_197 = (_zz_when_ArraySlice_l165_197 <= selectWriteFifo);
  assign when_ArraySlice_l166_197 = (_zz_when_ArraySlice_l166_197 <= _zz_when_ArraySlice_l166_197_2);
  assign _zz_when_ArraySlice_l112_197 = (wReg % _zz__zz_when_ArraySlice_l112_197);
  assign when_ArraySlice_l112_197 = (_zz_when_ArraySlice_l112_197 != 6'h0);
  assign when_ArraySlice_l113_197 = (7'h40 <= _zz_when_ArraySlice_l113_197);
  always @(*) begin
    if(when_ArraySlice_l112_197) begin
      if(when_ArraySlice_l113_197) begin
        _zz_when_ArraySlice_l173_197 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_197 = (_zz__zz_when_ArraySlice_l173_197 - _zz__zz_when_ArraySlice_l173_197_3);
      end
    end else begin
      if(when_ArraySlice_l118_197) begin
        _zz_when_ArraySlice_l173_197 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_197 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_197 = (_zz_when_ArraySlice_l118_197 <= wReg);
  assign when_ArraySlice_l173_197 = (_zz_when_ArraySlice_l173_197_1 <= _zz_when_ArraySlice_l173_197_3);
  assign when_ArraySlice_l165_198 = (_zz_when_ArraySlice_l165_198 <= selectWriteFifo);
  assign when_ArraySlice_l166_198 = (_zz_when_ArraySlice_l166_198 <= _zz_when_ArraySlice_l166_198_2);
  assign _zz_when_ArraySlice_l112_198 = (wReg % _zz__zz_when_ArraySlice_l112_198);
  assign when_ArraySlice_l112_198 = (_zz_when_ArraySlice_l112_198 != 6'h0);
  assign when_ArraySlice_l113_198 = (7'h40 <= _zz_when_ArraySlice_l113_198);
  always @(*) begin
    if(when_ArraySlice_l112_198) begin
      if(when_ArraySlice_l113_198) begin
        _zz_when_ArraySlice_l173_198 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_198 = (_zz__zz_when_ArraySlice_l173_198 - _zz__zz_when_ArraySlice_l173_198_3);
      end
    end else begin
      if(when_ArraySlice_l118_198) begin
        _zz_when_ArraySlice_l173_198 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_198 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_198 = (_zz_when_ArraySlice_l118_198 <= wReg);
  assign when_ArraySlice_l173_198 = (_zz_when_ArraySlice_l173_198_1 <= _zz_when_ArraySlice_l173_198_3);
  assign when_ArraySlice_l165_199 = (_zz_when_ArraySlice_l165_199 <= selectWriteFifo);
  assign when_ArraySlice_l166_199 = (_zz_when_ArraySlice_l166_199 <= _zz_when_ArraySlice_l166_199_2);
  assign _zz_when_ArraySlice_l112_199 = (wReg % _zz__zz_when_ArraySlice_l112_199);
  assign when_ArraySlice_l112_199 = (_zz_when_ArraySlice_l112_199 != 6'h0);
  assign when_ArraySlice_l113_199 = (7'h40 <= _zz_when_ArraySlice_l113_199);
  always @(*) begin
    if(when_ArraySlice_l112_199) begin
      if(when_ArraySlice_l113_199) begin
        _zz_when_ArraySlice_l173_199 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_199 = (_zz__zz_when_ArraySlice_l173_199 - _zz__zz_when_ArraySlice_l173_199_3);
      end
    end else begin
      if(when_ArraySlice_l118_199) begin
        _zz_when_ArraySlice_l173_199 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_199 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_199 = (_zz_when_ArraySlice_l118_199 <= wReg);
  assign when_ArraySlice_l173_199 = (_zz_when_ArraySlice_l173_199_1 <= _zz_when_ArraySlice_l173_199_3);
  assign when_ArraySlice_l444_7 = (! ((((((_zz_when_ArraySlice_l444_7 && _zz_when_ArraySlice_l444_7_1) && (holdReadOp_4 == _zz_when_ArraySlice_l444_7_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l444_7_3 && _zz_when_ArraySlice_l444_7_4) && (debug_4_24 == _zz_when_ArraySlice_l444_7_5)) && (debug_5_24 == 1'b1)) && (debug_6_24 == 1'b1)) && (debug_7_24 == 1'b1))));
  assign outputStreamArrayData_7_fire_5 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l448_7 = ((_zz_when_ArraySlice_l448_7 == 13'h0) && outputStreamArrayData_7_fire_5);
  assign when_ArraySlice_l434_7 = (allowPadding_7 && (wReg <= _zz_when_ArraySlice_l434_7));
  assign outputStreamArrayData_7_fire_6 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l455_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l455_7);
  always @(*) begin
    debug_0_25 = 1'b0;
    if(when_ArraySlice_l165_200) begin
      if(when_ArraySlice_l166_200) begin
        debug_0_25 = 1'b1;
      end else begin
        debug_0_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_200) begin
        debug_0_25 = 1'b1;
      end else begin
        debug_0_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_25 = 1'b0;
    if(when_ArraySlice_l165_201) begin
      if(when_ArraySlice_l166_201) begin
        debug_1_25 = 1'b1;
      end else begin
        debug_1_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_201) begin
        debug_1_25 = 1'b1;
      end else begin
        debug_1_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_25 = 1'b0;
    if(when_ArraySlice_l165_202) begin
      if(when_ArraySlice_l166_202) begin
        debug_2_25 = 1'b1;
      end else begin
        debug_2_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_202) begin
        debug_2_25 = 1'b1;
      end else begin
        debug_2_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_25 = 1'b0;
    if(when_ArraySlice_l165_203) begin
      if(when_ArraySlice_l166_203) begin
        debug_3_25 = 1'b1;
      end else begin
        debug_3_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_203) begin
        debug_3_25 = 1'b1;
      end else begin
        debug_3_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_25 = 1'b0;
    if(when_ArraySlice_l165_204) begin
      if(when_ArraySlice_l166_204) begin
        debug_4_25 = 1'b1;
      end else begin
        debug_4_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_204) begin
        debug_4_25 = 1'b1;
      end else begin
        debug_4_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_25 = 1'b0;
    if(when_ArraySlice_l165_205) begin
      if(when_ArraySlice_l166_205) begin
        debug_5_25 = 1'b1;
      end else begin
        debug_5_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_205) begin
        debug_5_25 = 1'b1;
      end else begin
        debug_5_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_25 = 1'b0;
    if(when_ArraySlice_l165_206) begin
      if(when_ArraySlice_l166_206) begin
        debug_6_25 = 1'b1;
      end else begin
        debug_6_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_206) begin
        debug_6_25 = 1'b1;
      end else begin
        debug_6_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_25 = 1'b0;
    if(when_ArraySlice_l165_207) begin
      if(when_ArraySlice_l166_207) begin
        debug_7_25 = 1'b1;
      end else begin
        debug_7_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_207) begin
        debug_7_25 = 1'b1;
      end else begin
        debug_7_25 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_200 = (_zz_when_ArraySlice_l165_200 <= selectWriteFifo);
  assign when_ArraySlice_l166_200 = (_zz_when_ArraySlice_l166_200 <= _zz_when_ArraySlice_l166_200_1);
  assign _zz_when_ArraySlice_l112_200 = (wReg % _zz__zz_when_ArraySlice_l112_200);
  assign when_ArraySlice_l112_200 = (_zz_when_ArraySlice_l112_200 != 6'h0);
  assign when_ArraySlice_l113_200 = (7'h40 <= _zz_when_ArraySlice_l113_200);
  always @(*) begin
    if(when_ArraySlice_l112_200) begin
      if(when_ArraySlice_l113_200) begin
        _zz_when_ArraySlice_l173_200 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_200 = (_zz__zz_when_ArraySlice_l173_200 - _zz__zz_when_ArraySlice_l173_200_3);
      end
    end else begin
      if(when_ArraySlice_l118_200) begin
        _zz_when_ArraySlice_l173_200 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_200 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_200 = (_zz_when_ArraySlice_l118_200 <= wReg);
  assign when_ArraySlice_l173_200 = (_zz_when_ArraySlice_l173_200_1 <= _zz_when_ArraySlice_l173_200_2);
  assign when_ArraySlice_l165_201 = (_zz_when_ArraySlice_l165_201 <= selectWriteFifo);
  assign when_ArraySlice_l166_201 = (_zz_when_ArraySlice_l166_201 <= _zz_when_ArraySlice_l166_201_1);
  assign _zz_when_ArraySlice_l112_201 = (wReg % _zz__zz_when_ArraySlice_l112_201);
  assign when_ArraySlice_l112_201 = (_zz_when_ArraySlice_l112_201 != 6'h0);
  assign when_ArraySlice_l113_201 = (7'h40 <= _zz_when_ArraySlice_l113_201);
  always @(*) begin
    if(when_ArraySlice_l112_201) begin
      if(when_ArraySlice_l113_201) begin
        _zz_when_ArraySlice_l173_201 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_201 = (_zz__zz_when_ArraySlice_l173_201 - _zz__zz_when_ArraySlice_l173_201_3);
      end
    end else begin
      if(when_ArraySlice_l118_201) begin
        _zz_when_ArraySlice_l173_201 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_201 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_201 = (_zz_when_ArraySlice_l118_201 <= wReg);
  assign when_ArraySlice_l173_201 = (_zz_when_ArraySlice_l173_201_1 <= _zz_when_ArraySlice_l173_201_3);
  assign when_ArraySlice_l165_202 = (_zz_when_ArraySlice_l165_202 <= selectWriteFifo);
  assign when_ArraySlice_l166_202 = (_zz_when_ArraySlice_l166_202 <= _zz_when_ArraySlice_l166_202_1);
  assign _zz_when_ArraySlice_l112_202 = (wReg % _zz__zz_when_ArraySlice_l112_202);
  assign when_ArraySlice_l112_202 = (_zz_when_ArraySlice_l112_202 != 6'h0);
  assign when_ArraySlice_l113_202 = (7'h40 <= _zz_when_ArraySlice_l113_202);
  always @(*) begin
    if(when_ArraySlice_l112_202) begin
      if(when_ArraySlice_l113_202) begin
        _zz_when_ArraySlice_l173_202 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_202 = (_zz__zz_when_ArraySlice_l173_202 - _zz__zz_when_ArraySlice_l173_202_3);
      end
    end else begin
      if(when_ArraySlice_l118_202) begin
        _zz_when_ArraySlice_l173_202 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_202 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_202 = (_zz_when_ArraySlice_l118_202 <= wReg);
  assign when_ArraySlice_l173_202 = (_zz_when_ArraySlice_l173_202_1 <= _zz_when_ArraySlice_l173_202_3);
  assign when_ArraySlice_l165_203 = (_zz_when_ArraySlice_l165_203 <= selectWriteFifo);
  assign when_ArraySlice_l166_203 = (_zz_when_ArraySlice_l166_203 <= _zz_when_ArraySlice_l166_203_1);
  assign _zz_when_ArraySlice_l112_203 = (wReg % _zz__zz_when_ArraySlice_l112_203);
  assign when_ArraySlice_l112_203 = (_zz_when_ArraySlice_l112_203 != 6'h0);
  assign when_ArraySlice_l113_203 = (7'h40 <= _zz_when_ArraySlice_l113_203);
  always @(*) begin
    if(when_ArraySlice_l112_203) begin
      if(when_ArraySlice_l113_203) begin
        _zz_when_ArraySlice_l173_203 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_203 = (_zz__zz_when_ArraySlice_l173_203 - _zz__zz_when_ArraySlice_l173_203_3);
      end
    end else begin
      if(when_ArraySlice_l118_203) begin
        _zz_when_ArraySlice_l173_203 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_203 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_203 = (_zz_when_ArraySlice_l118_203 <= wReg);
  assign when_ArraySlice_l173_203 = (_zz_when_ArraySlice_l173_203_1 <= _zz_when_ArraySlice_l173_203_3);
  assign when_ArraySlice_l165_204 = (_zz_when_ArraySlice_l165_204 <= selectWriteFifo);
  assign when_ArraySlice_l166_204 = (_zz_when_ArraySlice_l166_204 <= _zz_when_ArraySlice_l166_204_1);
  assign _zz_when_ArraySlice_l112_204 = (wReg % _zz__zz_when_ArraySlice_l112_204);
  assign when_ArraySlice_l112_204 = (_zz_when_ArraySlice_l112_204 != 6'h0);
  assign when_ArraySlice_l113_204 = (7'h40 <= _zz_when_ArraySlice_l113_204);
  always @(*) begin
    if(when_ArraySlice_l112_204) begin
      if(when_ArraySlice_l113_204) begin
        _zz_when_ArraySlice_l173_204 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_204 = (_zz__zz_when_ArraySlice_l173_204 - _zz__zz_when_ArraySlice_l173_204_3);
      end
    end else begin
      if(when_ArraySlice_l118_204) begin
        _zz_when_ArraySlice_l173_204 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_204 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_204 = (_zz_when_ArraySlice_l118_204 <= wReg);
  assign when_ArraySlice_l173_204 = (_zz_when_ArraySlice_l173_204_1 <= _zz_when_ArraySlice_l173_204_3);
  assign when_ArraySlice_l165_205 = (_zz_when_ArraySlice_l165_205 <= selectWriteFifo);
  assign when_ArraySlice_l166_205 = (_zz_when_ArraySlice_l166_205 <= _zz_when_ArraySlice_l166_205_2);
  assign _zz_when_ArraySlice_l112_205 = (wReg % _zz__zz_when_ArraySlice_l112_205);
  assign when_ArraySlice_l112_205 = (_zz_when_ArraySlice_l112_205 != 6'h0);
  assign when_ArraySlice_l113_205 = (7'h40 <= _zz_when_ArraySlice_l113_205);
  always @(*) begin
    if(when_ArraySlice_l112_205) begin
      if(when_ArraySlice_l113_205) begin
        _zz_when_ArraySlice_l173_205 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_205 = (_zz__zz_when_ArraySlice_l173_205 - _zz__zz_when_ArraySlice_l173_205_3);
      end
    end else begin
      if(when_ArraySlice_l118_205) begin
        _zz_when_ArraySlice_l173_205 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_205 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_205 = (_zz_when_ArraySlice_l118_205 <= wReg);
  assign when_ArraySlice_l173_205 = (_zz_when_ArraySlice_l173_205_1 <= _zz_when_ArraySlice_l173_205_3);
  assign when_ArraySlice_l165_206 = (_zz_when_ArraySlice_l165_206 <= selectWriteFifo);
  assign when_ArraySlice_l166_206 = (_zz_when_ArraySlice_l166_206 <= _zz_when_ArraySlice_l166_206_2);
  assign _zz_when_ArraySlice_l112_206 = (wReg % _zz__zz_when_ArraySlice_l112_206);
  assign when_ArraySlice_l112_206 = (_zz_when_ArraySlice_l112_206 != 6'h0);
  assign when_ArraySlice_l113_206 = (7'h40 <= _zz_when_ArraySlice_l113_206);
  always @(*) begin
    if(when_ArraySlice_l112_206) begin
      if(when_ArraySlice_l113_206) begin
        _zz_when_ArraySlice_l173_206 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_206 = (_zz__zz_when_ArraySlice_l173_206 - _zz__zz_when_ArraySlice_l173_206_3);
      end
    end else begin
      if(when_ArraySlice_l118_206) begin
        _zz_when_ArraySlice_l173_206 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_206 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_206 = (_zz_when_ArraySlice_l118_206 <= wReg);
  assign when_ArraySlice_l173_206 = (_zz_when_ArraySlice_l173_206_1 <= _zz_when_ArraySlice_l173_206_3);
  assign when_ArraySlice_l165_207 = (_zz_when_ArraySlice_l165_207 <= selectWriteFifo);
  assign when_ArraySlice_l166_207 = (_zz_when_ArraySlice_l166_207 <= _zz_when_ArraySlice_l166_207_2);
  assign _zz_when_ArraySlice_l112_207 = (wReg % _zz__zz_when_ArraySlice_l112_207);
  assign when_ArraySlice_l112_207 = (_zz_when_ArraySlice_l112_207 != 6'h0);
  assign when_ArraySlice_l113_207 = (7'h40 <= _zz_when_ArraySlice_l113_207);
  always @(*) begin
    if(when_ArraySlice_l112_207) begin
      if(when_ArraySlice_l113_207) begin
        _zz_when_ArraySlice_l173_207 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_207 = (_zz__zz_when_ArraySlice_l173_207 - _zz__zz_when_ArraySlice_l173_207_3);
      end
    end else begin
      if(when_ArraySlice_l118_207) begin
        _zz_when_ArraySlice_l173_207 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_207 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_207 = (_zz_when_ArraySlice_l118_207 <= wReg);
  assign when_ArraySlice_l173_207 = (_zz_when_ArraySlice_l173_207_1 <= _zz_when_ArraySlice_l173_207_3);
  assign when_ArraySlice_l465 = ((((((_zz_when_ArraySlice_l465 && _zz_when_ArraySlice_l465_1) && (holdReadOp_4 == _zz_when_ArraySlice_l465_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l465_3 && _zz_when_ArraySlice_l465_4) && (debug_4_25 == _zz_when_ArraySlice_l465_5)) && (debug_5_25 == 1'b1)) && (debug_6_25 == 1'b1)) && (debug_7_25 == 1'b1)));
  assign when_ArraySlice_l468 = (! allowPadding_0);
  assign when_ArraySlice_l468_1 = (! allowPadding_1);
  assign when_ArraySlice_l468_2 = (! allowPadding_2);
  assign when_ArraySlice_l468_3 = (! allowPadding_3);
  assign when_ArraySlice_l468_4 = (! allowPadding_4);
  assign when_ArraySlice_l468_5 = (! allowPadding_5);
  assign when_ArraySlice_l468_6 = (! allowPadding_6);
  assign when_ArraySlice_l468_7 = (! allowPadding_7);
  assign when_ArraySlice_l240 = (_zz_when_ArraySlice_l240 < wReg);
  assign when_ArraySlice_l241 = ((! holdReadOp_0) && (_zz_when_ArraySlice_l241 != 7'h0));
  assign _zz_outputStreamArrayData_0_valid_1 = (selectReadFifo_0 + _zz__zz_outputStreamArrayData_0_valid_1_1);
  assign _zz_11 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_0_valid_1);
  assign _zz_io_pop_ready_8 = outputStreamArrayData_0_ready;
  assign when_ArraySlice_l246 = (! holdReadOp_0);
  assign outputStreamArrayData_0_fire_7 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l247 = ((_zz_when_ArraySlice_l247 < _zz_when_ArraySlice_l247_2) && outputStreamArrayData_0_fire_7);
  assign when_ArraySlice_l248 = (handshakeTimes_0_value == _zz_when_ArraySlice_l248);
  assign when_ArraySlice_l251 = (_zz_when_ArraySlice_l251 == 13'h0);
  assign outputStreamArrayData_0_fire_8 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l256 = ((_zz_when_ArraySlice_l256 == _zz_when_ArraySlice_l256_4) && outputStreamArrayData_0_fire_8);
  assign when_ArraySlice_l257 = (handshakeTimes_0_value == _zz_when_ArraySlice_l257);
  assign _zz_when_ArraySlice_l94_24 = (hReg % _zz__zz_when_ArraySlice_l94_24);
  assign when_ArraySlice_l94_24 = (_zz_when_ArraySlice_l94_24 != 6'h0);
  assign when_ArraySlice_l95_24 = (7'h40 <= _zz_when_ArraySlice_l95_24);
  always @(*) begin
    if(when_ArraySlice_l94_24) begin
      if(when_ArraySlice_l95_24) begin
        _zz_when_ArraySlice_l259 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259 = (_zz__zz_when_ArraySlice_l259 - _zz__zz_when_ArraySlice_l259_3);
      end
    end else begin
      if(when_ArraySlice_l99_24) begin
        _zz_when_ArraySlice_l259 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_24 = (_zz_when_ArraySlice_l99_24 <= hReg);
  assign when_ArraySlice_l259 = (_zz_when_ArraySlice_l259_8 < _zz_when_ArraySlice_l259_11);
  always @(*) begin
    debug_0_26 = 1'b0;
    if(when_ArraySlice_l165_208) begin
      if(when_ArraySlice_l166_208) begin
        debug_0_26 = 1'b1;
      end else begin
        debug_0_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_208) begin
        debug_0_26 = 1'b1;
      end else begin
        debug_0_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_26 = 1'b0;
    if(when_ArraySlice_l165_209) begin
      if(when_ArraySlice_l166_209) begin
        debug_1_26 = 1'b1;
      end else begin
        debug_1_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_209) begin
        debug_1_26 = 1'b1;
      end else begin
        debug_1_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_26 = 1'b0;
    if(when_ArraySlice_l165_210) begin
      if(when_ArraySlice_l166_210) begin
        debug_2_26 = 1'b1;
      end else begin
        debug_2_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_210) begin
        debug_2_26 = 1'b1;
      end else begin
        debug_2_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_26 = 1'b0;
    if(when_ArraySlice_l165_211) begin
      if(when_ArraySlice_l166_211) begin
        debug_3_26 = 1'b1;
      end else begin
        debug_3_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_211) begin
        debug_3_26 = 1'b1;
      end else begin
        debug_3_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_26 = 1'b0;
    if(when_ArraySlice_l165_212) begin
      if(when_ArraySlice_l166_212) begin
        debug_4_26 = 1'b1;
      end else begin
        debug_4_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_212) begin
        debug_4_26 = 1'b1;
      end else begin
        debug_4_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_26 = 1'b0;
    if(when_ArraySlice_l165_213) begin
      if(when_ArraySlice_l166_213) begin
        debug_5_26 = 1'b1;
      end else begin
        debug_5_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_213) begin
        debug_5_26 = 1'b1;
      end else begin
        debug_5_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_26 = 1'b0;
    if(when_ArraySlice_l165_214) begin
      if(when_ArraySlice_l166_214) begin
        debug_6_26 = 1'b1;
      end else begin
        debug_6_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_214) begin
        debug_6_26 = 1'b1;
      end else begin
        debug_6_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_26 = 1'b0;
    if(when_ArraySlice_l165_215) begin
      if(when_ArraySlice_l166_215) begin
        debug_7_26 = 1'b1;
      end else begin
        debug_7_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_215) begin
        debug_7_26 = 1'b1;
      end else begin
        debug_7_26 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_208 = (_zz_when_ArraySlice_l165_208 <= selectWriteFifo);
  assign when_ArraySlice_l166_208 = (_zz_when_ArraySlice_l166_208 <= _zz_when_ArraySlice_l166_208_1);
  assign _zz_when_ArraySlice_l112_208 = (wReg % _zz__zz_when_ArraySlice_l112_208);
  assign when_ArraySlice_l112_208 = (_zz_when_ArraySlice_l112_208 != 6'h0);
  assign when_ArraySlice_l113_208 = (7'h40 <= _zz_when_ArraySlice_l113_208);
  always @(*) begin
    if(when_ArraySlice_l112_208) begin
      if(when_ArraySlice_l113_208) begin
        _zz_when_ArraySlice_l173_208 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_208 = (_zz__zz_when_ArraySlice_l173_208 - _zz__zz_when_ArraySlice_l173_208_3);
      end
    end else begin
      if(when_ArraySlice_l118_208) begin
        _zz_when_ArraySlice_l173_208 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_208 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_208 = (_zz_when_ArraySlice_l118_208 <= wReg);
  assign when_ArraySlice_l173_208 = (_zz_when_ArraySlice_l173_208_1 <= _zz_when_ArraySlice_l173_208_2);
  assign when_ArraySlice_l165_209 = (_zz_when_ArraySlice_l165_209 <= selectWriteFifo);
  assign when_ArraySlice_l166_209 = (_zz_when_ArraySlice_l166_209 <= _zz_when_ArraySlice_l166_209_1);
  assign _zz_when_ArraySlice_l112_209 = (wReg % _zz__zz_when_ArraySlice_l112_209);
  assign when_ArraySlice_l112_209 = (_zz_when_ArraySlice_l112_209 != 6'h0);
  assign when_ArraySlice_l113_209 = (7'h40 <= _zz_when_ArraySlice_l113_209);
  always @(*) begin
    if(when_ArraySlice_l112_209) begin
      if(when_ArraySlice_l113_209) begin
        _zz_when_ArraySlice_l173_209 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_209 = (_zz__zz_when_ArraySlice_l173_209 - _zz__zz_when_ArraySlice_l173_209_3);
      end
    end else begin
      if(when_ArraySlice_l118_209) begin
        _zz_when_ArraySlice_l173_209 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_209 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_209 = (_zz_when_ArraySlice_l118_209 <= wReg);
  assign when_ArraySlice_l173_209 = (_zz_when_ArraySlice_l173_209_1 <= _zz_when_ArraySlice_l173_209_3);
  assign when_ArraySlice_l165_210 = (_zz_when_ArraySlice_l165_210 <= selectWriteFifo);
  assign when_ArraySlice_l166_210 = (_zz_when_ArraySlice_l166_210 <= _zz_when_ArraySlice_l166_210_1);
  assign _zz_when_ArraySlice_l112_210 = (wReg % _zz__zz_when_ArraySlice_l112_210);
  assign when_ArraySlice_l112_210 = (_zz_when_ArraySlice_l112_210 != 6'h0);
  assign when_ArraySlice_l113_210 = (7'h40 <= _zz_when_ArraySlice_l113_210);
  always @(*) begin
    if(when_ArraySlice_l112_210) begin
      if(when_ArraySlice_l113_210) begin
        _zz_when_ArraySlice_l173_210 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_210 = (_zz__zz_when_ArraySlice_l173_210 - _zz__zz_when_ArraySlice_l173_210_3);
      end
    end else begin
      if(when_ArraySlice_l118_210) begin
        _zz_when_ArraySlice_l173_210 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_210 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_210 = (_zz_when_ArraySlice_l118_210 <= wReg);
  assign when_ArraySlice_l173_210 = (_zz_when_ArraySlice_l173_210_1 <= _zz_when_ArraySlice_l173_210_3);
  assign when_ArraySlice_l165_211 = (_zz_when_ArraySlice_l165_211 <= selectWriteFifo);
  assign when_ArraySlice_l166_211 = (_zz_when_ArraySlice_l166_211 <= _zz_when_ArraySlice_l166_211_1);
  assign _zz_when_ArraySlice_l112_211 = (wReg % _zz__zz_when_ArraySlice_l112_211);
  assign when_ArraySlice_l112_211 = (_zz_when_ArraySlice_l112_211 != 6'h0);
  assign when_ArraySlice_l113_211 = (7'h40 <= _zz_when_ArraySlice_l113_211);
  always @(*) begin
    if(when_ArraySlice_l112_211) begin
      if(when_ArraySlice_l113_211) begin
        _zz_when_ArraySlice_l173_211 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_211 = (_zz__zz_when_ArraySlice_l173_211 - _zz__zz_when_ArraySlice_l173_211_3);
      end
    end else begin
      if(when_ArraySlice_l118_211) begin
        _zz_when_ArraySlice_l173_211 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_211 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_211 = (_zz_when_ArraySlice_l118_211 <= wReg);
  assign when_ArraySlice_l173_211 = (_zz_when_ArraySlice_l173_211_1 <= _zz_when_ArraySlice_l173_211_3);
  assign when_ArraySlice_l165_212 = (_zz_when_ArraySlice_l165_212 <= selectWriteFifo);
  assign when_ArraySlice_l166_212 = (_zz_when_ArraySlice_l166_212 <= _zz_when_ArraySlice_l166_212_1);
  assign _zz_when_ArraySlice_l112_212 = (wReg % _zz__zz_when_ArraySlice_l112_212);
  assign when_ArraySlice_l112_212 = (_zz_when_ArraySlice_l112_212 != 6'h0);
  assign when_ArraySlice_l113_212 = (7'h40 <= _zz_when_ArraySlice_l113_212);
  always @(*) begin
    if(when_ArraySlice_l112_212) begin
      if(when_ArraySlice_l113_212) begin
        _zz_when_ArraySlice_l173_212 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_212 = (_zz__zz_when_ArraySlice_l173_212 - _zz__zz_when_ArraySlice_l173_212_3);
      end
    end else begin
      if(when_ArraySlice_l118_212) begin
        _zz_when_ArraySlice_l173_212 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_212 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_212 = (_zz_when_ArraySlice_l118_212 <= wReg);
  assign when_ArraySlice_l173_212 = (_zz_when_ArraySlice_l173_212_1 <= _zz_when_ArraySlice_l173_212_3);
  assign when_ArraySlice_l165_213 = (_zz_when_ArraySlice_l165_213 <= selectWriteFifo);
  assign when_ArraySlice_l166_213 = (_zz_when_ArraySlice_l166_213 <= _zz_when_ArraySlice_l166_213_2);
  assign _zz_when_ArraySlice_l112_213 = (wReg % _zz__zz_when_ArraySlice_l112_213);
  assign when_ArraySlice_l112_213 = (_zz_when_ArraySlice_l112_213 != 6'h0);
  assign when_ArraySlice_l113_213 = (7'h40 <= _zz_when_ArraySlice_l113_213);
  always @(*) begin
    if(when_ArraySlice_l112_213) begin
      if(when_ArraySlice_l113_213) begin
        _zz_when_ArraySlice_l173_213 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_213 = (_zz__zz_when_ArraySlice_l173_213 - _zz__zz_when_ArraySlice_l173_213_3);
      end
    end else begin
      if(when_ArraySlice_l118_213) begin
        _zz_when_ArraySlice_l173_213 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_213 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_213 = (_zz_when_ArraySlice_l118_213 <= wReg);
  assign when_ArraySlice_l173_213 = (_zz_when_ArraySlice_l173_213_1 <= _zz_when_ArraySlice_l173_213_3);
  assign when_ArraySlice_l165_214 = (_zz_when_ArraySlice_l165_214 <= selectWriteFifo);
  assign when_ArraySlice_l166_214 = (_zz_when_ArraySlice_l166_214 <= _zz_when_ArraySlice_l166_214_2);
  assign _zz_when_ArraySlice_l112_214 = (wReg % _zz__zz_when_ArraySlice_l112_214);
  assign when_ArraySlice_l112_214 = (_zz_when_ArraySlice_l112_214 != 6'h0);
  assign when_ArraySlice_l113_214 = (7'h40 <= _zz_when_ArraySlice_l113_214);
  always @(*) begin
    if(when_ArraySlice_l112_214) begin
      if(when_ArraySlice_l113_214) begin
        _zz_when_ArraySlice_l173_214 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_214 = (_zz__zz_when_ArraySlice_l173_214 - _zz__zz_when_ArraySlice_l173_214_3);
      end
    end else begin
      if(when_ArraySlice_l118_214) begin
        _zz_when_ArraySlice_l173_214 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_214 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_214 = (_zz_when_ArraySlice_l118_214 <= wReg);
  assign when_ArraySlice_l173_214 = (_zz_when_ArraySlice_l173_214_1 <= _zz_when_ArraySlice_l173_214_3);
  assign when_ArraySlice_l165_215 = (_zz_when_ArraySlice_l165_215 <= selectWriteFifo);
  assign when_ArraySlice_l166_215 = (_zz_when_ArraySlice_l166_215 <= _zz_when_ArraySlice_l166_215_2);
  assign _zz_when_ArraySlice_l112_215 = (wReg % _zz__zz_when_ArraySlice_l112_215);
  assign when_ArraySlice_l112_215 = (_zz_when_ArraySlice_l112_215 != 6'h0);
  assign when_ArraySlice_l113_215 = (7'h40 <= _zz_when_ArraySlice_l113_215);
  always @(*) begin
    if(when_ArraySlice_l112_215) begin
      if(when_ArraySlice_l113_215) begin
        _zz_when_ArraySlice_l173_215 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_215 = (_zz__zz_when_ArraySlice_l173_215 - _zz__zz_when_ArraySlice_l173_215_3);
      end
    end else begin
      if(when_ArraySlice_l118_215) begin
        _zz_when_ArraySlice_l173_215 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_215 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_215 = (_zz_when_ArraySlice_l118_215 <= wReg);
  assign when_ArraySlice_l173_215 = (_zz_when_ArraySlice_l173_215_1 <= _zz_when_ArraySlice_l173_215_3);
  assign when_ArraySlice_l265 = (! ((((((_zz_when_ArraySlice_l265 && _zz_when_ArraySlice_l265_1) && (holdReadOp_4 == _zz_when_ArraySlice_l265_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l265_3 && _zz_when_ArraySlice_l265_4) && (debug_4_26 == _zz_when_ArraySlice_l265_5)) && (debug_5_26 == 1'b1)) && (debug_6_26 == 1'b1)) && (debug_7_26 == 1'b1))));
  assign when_ArraySlice_l268 = (wReg <= _zz_when_ArraySlice_l268);
  assign when_ArraySlice_l272 = (_zz_when_ArraySlice_l272 == 13'h0);
  assign when_ArraySlice_l276 = (_zz_when_ArraySlice_l276 == 7'h0);
  assign outputStreamArrayData_0_fire_9 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l277 = ((handshakeTimes_0_value == _zz_when_ArraySlice_l277) && outputStreamArrayData_0_fire_9);
  assign _zz_when_ArraySlice_l94_25 = (hReg % _zz__zz_when_ArraySlice_l94_25);
  assign when_ArraySlice_l94_25 = (_zz_when_ArraySlice_l94_25 != 6'h0);
  assign when_ArraySlice_l95_25 = (7'h40 <= _zz_when_ArraySlice_l95_25);
  always @(*) begin
    if(when_ArraySlice_l94_25) begin
      if(when_ArraySlice_l95_25) begin
        _zz_when_ArraySlice_l279 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279 = (_zz__zz_when_ArraySlice_l279 - _zz__zz_when_ArraySlice_l279_3);
      end
    end else begin
      if(when_ArraySlice_l99_25) begin
        _zz_when_ArraySlice_l279 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_25 = (_zz_when_ArraySlice_l99_25 <= hReg);
  assign when_ArraySlice_l279 = (_zz_when_ArraySlice_l279_8 < _zz_when_ArraySlice_l279_11);
  always @(*) begin
    debug_0_27 = 1'b0;
    if(when_ArraySlice_l165_216) begin
      if(when_ArraySlice_l166_216) begin
        debug_0_27 = 1'b1;
      end else begin
        debug_0_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_216) begin
        debug_0_27 = 1'b1;
      end else begin
        debug_0_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_27 = 1'b0;
    if(when_ArraySlice_l165_217) begin
      if(when_ArraySlice_l166_217) begin
        debug_1_27 = 1'b1;
      end else begin
        debug_1_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_217) begin
        debug_1_27 = 1'b1;
      end else begin
        debug_1_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_27 = 1'b0;
    if(when_ArraySlice_l165_218) begin
      if(when_ArraySlice_l166_218) begin
        debug_2_27 = 1'b1;
      end else begin
        debug_2_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_218) begin
        debug_2_27 = 1'b1;
      end else begin
        debug_2_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_27 = 1'b0;
    if(when_ArraySlice_l165_219) begin
      if(when_ArraySlice_l166_219) begin
        debug_3_27 = 1'b1;
      end else begin
        debug_3_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_219) begin
        debug_3_27 = 1'b1;
      end else begin
        debug_3_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_27 = 1'b0;
    if(when_ArraySlice_l165_220) begin
      if(when_ArraySlice_l166_220) begin
        debug_4_27 = 1'b1;
      end else begin
        debug_4_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_220) begin
        debug_4_27 = 1'b1;
      end else begin
        debug_4_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_27 = 1'b0;
    if(when_ArraySlice_l165_221) begin
      if(when_ArraySlice_l166_221) begin
        debug_5_27 = 1'b1;
      end else begin
        debug_5_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_221) begin
        debug_5_27 = 1'b1;
      end else begin
        debug_5_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_27 = 1'b0;
    if(when_ArraySlice_l165_222) begin
      if(when_ArraySlice_l166_222) begin
        debug_6_27 = 1'b1;
      end else begin
        debug_6_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_222) begin
        debug_6_27 = 1'b1;
      end else begin
        debug_6_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_27 = 1'b0;
    if(when_ArraySlice_l165_223) begin
      if(when_ArraySlice_l166_223) begin
        debug_7_27 = 1'b1;
      end else begin
        debug_7_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_223) begin
        debug_7_27 = 1'b1;
      end else begin
        debug_7_27 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_216 = (_zz_when_ArraySlice_l165_216 <= selectWriteFifo);
  assign when_ArraySlice_l166_216 = (_zz_when_ArraySlice_l166_216 <= _zz_when_ArraySlice_l166_216_1);
  assign _zz_when_ArraySlice_l112_216 = (wReg % _zz__zz_when_ArraySlice_l112_216);
  assign when_ArraySlice_l112_216 = (_zz_when_ArraySlice_l112_216 != 6'h0);
  assign when_ArraySlice_l113_216 = (7'h40 <= _zz_when_ArraySlice_l113_216);
  always @(*) begin
    if(when_ArraySlice_l112_216) begin
      if(when_ArraySlice_l113_216) begin
        _zz_when_ArraySlice_l173_216 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_216 = (_zz__zz_when_ArraySlice_l173_216 - _zz__zz_when_ArraySlice_l173_216_3);
      end
    end else begin
      if(when_ArraySlice_l118_216) begin
        _zz_when_ArraySlice_l173_216 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_216 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_216 = (_zz_when_ArraySlice_l118_216 <= wReg);
  assign when_ArraySlice_l173_216 = (_zz_when_ArraySlice_l173_216_1 <= _zz_when_ArraySlice_l173_216_2);
  assign when_ArraySlice_l165_217 = (_zz_when_ArraySlice_l165_217 <= selectWriteFifo);
  assign when_ArraySlice_l166_217 = (_zz_when_ArraySlice_l166_217 <= _zz_when_ArraySlice_l166_217_1);
  assign _zz_when_ArraySlice_l112_217 = (wReg % _zz__zz_when_ArraySlice_l112_217);
  assign when_ArraySlice_l112_217 = (_zz_when_ArraySlice_l112_217 != 6'h0);
  assign when_ArraySlice_l113_217 = (7'h40 <= _zz_when_ArraySlice_l113_217);
  always @(*) begin
    if(when_ArraySlice_l112_217) begin
      if(when_ArraySlice_l113_217) begin
        _zz_when_ArraySlice_l173_217 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_217 = (_zz__zz_when_ArraySlice_l173_217 - _zz__zz_when_ArraySlice_l173_217_3);
      end
    end else begin
      if(when_ArraySlice_l118_217) begin
        _zz_when_ArraySlice_l173_217 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_217 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_217 = (_zz_when_ArraySlice_l118_217 <= wReg);
  assign when_ArraySlice_l173_217 = (_zz_when_ArraySlice_l173_217_1 <= _zz_when_ArraySlice_l173_217_3);
  assign when_ArraySlice_l165_218 = (_zz_when_ArraySlice_l165_218 <= selectWriteFifo);
  assign when_ArraySlice_l166_218 = (_zz_when_ArraySlice_l166_218 <= _zz_when_ArraySlice_l166_218_1);
  assign _zz_when_ArraySlice_l112_218 = (wReg % _zz__zz_when_ArraySlice_l112_218);
  assign when_ArraySlice_l112_218 = (_zz_when_ArraySlice_l112_218 != 6'h0);
  assign when_ArraySlice_l113_218 = (7'h40 <= _zz_when_ArraySlice_l113_218);
  always @(*) begin
    if(when_ArraySlice_l112_218) begin
      if(when_ArraySlice_l113_218) begin
        _zz_when_ArraySlice_l173_218 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_218 = (_zz__zz_when_ArraySlice_l173_218 - _zz__zz_when_ArraySlice_l173_218_3);
      end
    end else begin
      if(when_ArraySlice_l118_218) begin
        _zz_when_ArraySlice_l173_218 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_218 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_218 = (_zz_when_ArraySlice_l118_218 <= wReg);
  assign when_ArraySlice_l173_218 = (_zz_when_ArraySlice_l173_218_1 <= _zz_when_ArraySlice_l173_218_3);
  assign when_ArraySlice_l165_219 = (_zz_when_ArraySlice_l165_219 <= selectWriteFifo);
  assign when_ArraySlice_l166_219 = (_zz_when_ArraySlice_l166_219 <= _zz_when_ArraySlice_l166_219_1);
  assign _zz_when_ArraySlice_l112_219 = (wReg % _zz__zz_when_ArraySlice_l112_219);
  assign when_ArraySlice_l112_219 = (_zz_when_ArraySlice_l112_219 != 6'h0);
  assign when_ArraySlice_l113_219 = (7'h40 <= _zz_when_ArraySlice_l113_219);
  always @(*) begin
    if(when_ArraySlice_l112_219) begin
      if(when_ArraySlice_l113_219) begin
        _zz_when_ArraySlice_l173_219 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_219 = (_zz__zz_when_ArraySlice_l173_219 - _zz__zz_when_ArraySlice_l173_219_3);
      end
    end else begin
      if(when_ArraySlice_l118_219) begin
        _zz_when_ArraySlice_l173_219 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_219 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_219 = (_zz_when_ArraySlice_l118_219 <= wReg);
  assign when_ArraySlice_l173_219 = (_zz_when_ArraySlice_l173_219_1 <= _zz_when_ArraySlice_l173_219_3);
  assign when_ArraySlice_l165_220 = (_zz_when_ArraySlice_l165_220 <= selectWriteFifo);
  assign when_ArraySlice_l166_220 = (_zz_when_ArraySlice_l166_220 <= _zz_when_ArraySlice_l166_220_1);
  assign _zz_when_ArraySlice_l112_220 = (wReg % _zz__zz_when_ArraySlice_l112_220);
  assign when_ArraySlice_l112_220 = (_zz_when_ArraySlice_l112_220 != 6'h0);
  assign when_ArraySlice_l113_220 = (7'h40 <= _zz_when_ArraySlice_l113_220);
  always @(*) begin
    if(when_ArraySlice_l112_220) begin
      if(when_ArraySlice_l113_220) begin
        _zz_when_ArraySlice_l173_220 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_220 = (_zz__zz_when_ArraySlice_l173_220 - _zz__zz_when_ArraySlice_l173_220_3);
      end
    end else begin
      if(when_ArraySlice_l118_220) begin
        _zz_when_ArraySlice_l173_220 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_220 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_220 = (_zz_when_ArraySlice_l118_220 <= wReg);
  assign when_ArraySlice_l173_220 = (_zz_when_ArraySlice_l173_220_1 <= _zz_when_ArraySlice_l173_220_3);
  assign when_ArraySlice_l165_221 = (_zz_when_ArraySlice_l165_221 <= selectWriteFifo);
  assign when_ArraySlice_l166_221 = (_zz_when_ArraySlice_l166_221 <= _zz_when_ArraySlice_l166_221_2);
  assign _zz_when_ArraySlice_l112_221 = (wReg % _zz__zz_when_ArraySlice_l112_221);
  assign when_ArraySlice_l112_221 = (_zz_when_ArraySlice_l112_221 != 6'h0);
  assign when_ArraySlice_l113_221 = (7'h40 <= _zz_when_ArraySlice_l113_221);
  always @(*) begin
    if(when_ArraySlice_l112_221) begin
      if(when_ArraySlice_l113_221) begin
        _zz_when_ArraySlice_l173_221 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_221 = (_zz__zz_when_ArraySlice_l173_221 - _zz__zz_when_ArraySlice_l173_221_3);
      end
    end else begin
      if(when_ArraySlice_l118_221) begin
        _zz_when_ArraySlice_l173_221 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_221 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_221 = (_zz_when_ArraySlice_l118_221 <= wReg);
  assign when_ArraySlice_l173_221 = (_zz_when_ArraySlice_l173_221_1 <= _zz_when_ArraySlice_l173_221_3);
  assign when_ArraySlice_l165_222 = (_zz_when_ArraySlice_l165_222 <= selectWriteFifo);
  assign when_ArraySlice_l166_222 = (_zz_when_ArraySlice_l166_222 <= _zz_when_ArraySlice_l166_222_2);
  assign _zz_when_ArraySlice_l112_222 = (wReg % _zz__zz_when_ArraySlice_l112_222);
  assign when_ArraySlice_l112_222 = (_zz_when_ArraySlice_l112_222 != 6'h0);
  assign when_ArraySlice_l113_222 = (7'h40 <= _zz_when_ArraySlice_l113_222);
  always @(*) begin
    if(when_ArraySlice_l112_222) begin
      if(when_ArraySlice_l113_222) begin
        _zz_when_ArraySlice_l173_222 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_222 = (_zz__zz_when_ArraySlice_l173_222 - _zz__zz_when_ArraySlice_l173_222_3);
      end
    end else begin
      if(when_ArraySlice_l118_222) begin
        _zz_when_ArraySlice_l173_222 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_222 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_222 = (_zz_when_ArraySlice_l118_222 <= wReg);
  assign when_ArraySlice_l173_222 = (_zz_when_ArraySlice_l173_222_1 <= _zz_when_ArraySlice_l173_222_3);
  assign when_ArraySlice_l165_223 = (_zz_when_ArraySlice_l165_223 <= selectWriteFifo);
  assign when_ArraySlice_l166_223 = (_zz_when_ArraySlice_l166_223 <= _zz_when_ArraySlice_l166_223_2);
  assign _zz_when_ArraySlice_l112_223 = (wReg % _zz__zz_when_ArraySlice_l112_223);
  assign when_ArraySlice_l112_223 = (_zz_when_ArraySlice_l112_223 != 6'h0);
  assign when_ArraySlice_l113_223 = (7'h40 <= _zz_when_ArraySlice_l113_223);
  always @(*) begin
    if(when_ArraySlice_l112_223) begin
      if(when_ArraySlice_l113_223) begin
        _zz_when_ArraySlice_l173_223 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_223 = (_zz__zz_when_ArraySlice_l173_223 - _zz__zz_when_ArraySlice_l173_223_3);
      end
    end else begin
      if(when_ArraySlice_l118_223) begin
        _zz_when_ArraySlice_l173_223 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_223 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_223 = (_zz_when_ArraySlice_l118_223 <= wReg);
  assign when_ArraySlice_l173_223 = (_zz_when_ArraySlice_l173_223_1 <= _zz_when_ArraySlice_l173_223_3);
  assign when_ArraySlice_l285 = (! ((((((_zz_when_ArraySlice_l285 && _zz_when_ArraySlice_l285_1) && (holdReadOp_4 == _zz_when_ArraySlice_l285_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l285_3 && _zz_when_ArraySlice_l285_4) && (debug_4_27 == _zz_when_ArraySlice_l285_5)) && (debug_5_27 == 1'b1)) && (debug_6_27 == 1'b1)) && (debug_7_27 == 1'b1))));
  assign when_ArraySlice_l288 = (wReg <= _zz_when_ArraySlice_l288);
  assign outputStreamArrayData_0_fire_10 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l292 = ((_zz_when_ArraySlice_l292 == 13'h0) && outputStreamArrayData_0_fire_10);
  assign outputStreamArrayData_0_fire_11 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l303 = ((handshakeTimes_0_value == _zz_when_ArraySlice_l303) && outputStreamArrayData_0_fire_11);
  assign _zz_when_ArraySlice_l94_26 = (hReg % _zz__zz_when_ArraySlice_l94_26);
  assign when_ArraySlice_l94_26 = (_zz_when_ArraySlice_l94_26 != 6'h0);
  assign when_ArraySlice_l95_26 = (7'h40 <= _zz_when_ArraySlice_l95_26);
  always @(*) begin
    if(when_ArraySlice_l94_26) begin
      if(when_ArraySlice_l95_26) begin
        _zz_when_ArraySlice_l304 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304 = (_zz__zz_when_ArraySlice_l304 - _zz__zz_when_ArraySlice_l304_3);
      end
    end else begin
      if(when_ArraySlice_l99_26) begin
        _zz_when_ArraySlice_l304 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_26 = (_zz_when_ArraySlice_l99_26 <= hReg);
  assign when_ArraySlice_l304 = (_zz_when_ArraySlice_l304_8 < _zz_when_ArraySlice_l304_11);
  always @(*) begin
    debug_0_28 = 1'b0;
    if(when_ArraySlice_l165_224) begin
      if(when_ArraySlice_l166_224) begin
        debug_0_28 = 1'b1;
      end else begin
        debug_0_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_224) begin
        debug_0_28 = 1'b1;
      end else begin
        debug_0_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_28 = 1'b0;
    if(when_ArraySlice_l165_225) begin
      if(when_ArraySlice_l166_225) begin
        debug_1_28 = 1'b1;
      end else begin
        debug_1_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_225) begin
        debug_1_28 = 1'b1;
      end else begin
        debug_1_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_28 = 1'b0;
    if(when_ArraySlice_l165_226) begin
      if(when_ArraySlice_l166_226) begin
        debug_2_28 = 1'b1;
      end else begin
        debug_2_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_226) begin
        debug_2_28 = 1'b1;
      end else begin
        debug_2_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_28 = 1'b0;
    if(when_ArraySlice_l165_227) begin
      if(when_ArraySlice_l166_227) begin
        debug_3_28 = 1'b1;
      end else begin
        debug_3_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_227) begin
        debug_3_28 = 1'b1;
      end else begin
        debug_3_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_28 = 1'b0;
    if(when_ArraySlice_l165_228) begin
      if(when_ArraySlice_l166_228) begin
        debug_4_28 = 1'b1;
      end else begin
        debug_4_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_228) begin
        debug_4_28 = 1'b1;
      end else begin
        debug_4_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_28 = 1'b0;
    if(when_ArraySlice_l165_229) begin
      if(when_ArraySlice_l166_229) begin
        debug_5_28 = 1'b1;
      end else begin
        debug_5_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_229) begin
        debug_5_28 = 1'b1;
      end else begin
        debug_5_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_28 = 1'b0;
    if(when_ArraySlice_l165_230) begin
      if(when_ArraySlice_l166_230) begin
        debug_6_28 = 1'b1;
      end else begin
        debug_6_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_230) begin
        debug_6_28 = 1'b1;
      end else begin
        debug_6_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_28 = 1'b0;
    if(when_ArraySlice_l165_231) begin
      if(when_ArraySlice_l166_231) begin
        debug_7_28 = 1'b1;
      end else begin
        debug_7_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_231) begin
        debug_7_28 = 1'b1;
      end else begin
        debug_7_28 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_224 = (_zz_when_ArraySlice_l165_224 <= selectWriteFifo);
  assign when_ArraySlice_l166_224 = (_zz_when_ArraySlice_l166_224 <= _zz_when_ArraySlice_l166_224_1);
  assign _zz_when_ArraySlice_l112_224 = (wReg % _zz__zz_when_ArraySlice_l112_224);
  assign when_ArraySlice_l112_224 = (_zz_when_ArraySlice_l112_224 != 6'h0);
  assign when_ArraySlice_l113_224 = (7'h40 <= _zz_when_ArraySlice_l113_224);
  always @(*) begin
    if(when_ArraySlice_l112_224) begin
      if(when_ArraySlice_l113_224) begin
        _zz_when_ArraySlice_l173_224 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_224 = (_zz__zz_when_ArraySlice_l173_224 - _zz__zz_when_ArraySlice_l173_224_3);
      end
    end else begin
      if(when_ArraySlice_l118_224) begin
        _zz_when_ArraySlice_l173_224 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_224 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_224 = (_zz_when_ArraySlice_l118_224 <= wReg);
  assign when_ArraySlice_l173_224 = (_zz_when_ArraySlice_l173_224_1 <= _zz_when_ArraySlice_l173_224_2);
  assign when_ArraySlice_l165_225 = (_zz_when_ArraySlice_l165_225 <= selectWriteFifo);
  assign when_ArraySlice_l166_225 = (_zz_when_ArraySlice_l166_225 <= _zz_when_ArraySlice_l166_225_1);
  assign _zz_when_ArraySlice_l112_225 = (wReg % _zz__zz_when_ArraySlice_l112_225);
  assign when_ArraySlice_l112_225 = (_zz_when_ArraySlice_l112_225 != 6'h0);
  assign when_ArraySlice_l113_225 = (7'h40 <= _zz_when_ArraySlice_l113_225);
  always @(*) begin
    if(when_ArraySlice_l112_225) begin
      if(when_ArraySlice_l113_225) begin
        _zz_when_ArraySlice_l173_225 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_225 = (_zz__zz_when_ArraySlice_l173_225 - _zz__zz_when_ArraySlice_l173_225_3);
      end
    end else begin
      if(when_ArraySlice_l118_225) begin
        _zz_when_ArraySlice_l173_225 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_225 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_225 = (_zz_when_ArraySlice_l118_225 <= wReg);
  assign when_ArraySlice_l173_225 = (_zz_when_ArraySlice_l173_225_1 <= _zz_when_ArraySlice_l173_225_3);
  assign when_ArraySlice_l165_226 = (_zz_when_ArraySlice_l165_226 <= selectWriteFifo);
  assign when_ArraySlice_l166_226 = (_zz_when_ArraySlice_l166_226 <= _zz_when_ArraySlice_l166_226_1);
  assign _zz_when_ArraySlice_l112_226 = (wReg % _zz__zz_when_ArraySlice_l112_226);
  assign when_ArraySlice_l112_226 = (_zz_when_ArraySlice_l112_226 != 6'h0);
  assign when_ArraySlice_l113_226 = (7'h40 <= _zz_when_ArraySlice_l113_226);
  always @(*) begin
    if(when_ArraySlice_l112_226) begin
      if(when_ArraySlice_l113_226) begin
        _zz_when_ArraySlice_l173_226 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_226 = (_zz__zz_when_ArraySlice_l173_226 - _zz__zz_when_ArraySlice_l173_226_3);
      end
    end else begin
      if(when_ArraySlice_l118_226) begin
        _zz_when_ArraySlice_l173_226 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_226 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_226 = (_zz_when_ArraySlice_l118_226 <= wReg);
  assign when_ArraySlice_l173_226 = (_zz_when_ArraySlice_l173_226_1 <= _zz_when_ArraySlice_l173_226_3);
  assign when_ArraySlice_l165_227 = (_zz_when_ArraySlice_l165_227 <= selectWriteFifo);
  assign when_ArraySlice_l166_227 = (_zz_when_ArraySlice_l166_227 <= _zz_when_ArraySlice_l166_227_1);
  assign _zz_when_ArraySlice_l112_227 = (wReg % _zz__zz_when_ArraySlice_l112_227);
  assign when_ArraySlice_l112_227 = (_zz_when_ArraySlice_l112_227 != 6'h0);
  assign when_ArraySlice_l113_227 = (7'h40 <= _zz_when_ArraySlice_l113_227);
  always @(*) begin
    if(when_ArraySlice_l112_227) begin
      if(when_ArraySlice_l113_227) begin
        _zz_when_ArraySlice_l173_227 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_227 = (_zz__zz_when_ArraySlice_l173_227 - _zz__zz_when_ArraySlice_l173_227_3);
      end
    end else begin
      if(when_ArraySlice_l118_227) begin
        _zz_when_ArraySlice_l173_227 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_227 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_227 = (_zz_when_ArraySlice_l118_227 <= wReg);
  assign when_ArraySlice_l173_227 = (_zz_when_ArraySlice_l173_227_1 <= _zz_when_ArraySlice_l173_227_3);
  assign when_ArraySlice_l165_228 = (_zz_when_ArraySlice_l165_228 <= selectWriteFifo);
  assign when_ArraySlice_l166_228 = (_zz_when_ArraySlice_l166_228 <= _zz_when_ArraySlice_l166_228_1);
  assign _zz_when_ArraySlice_l112_228 = (wReg % _zz__zz_when_ArraySlice_l112_228);
  assign when_ArraySlice_l112_228 = (_zz_when_ArraySlice_l112_228 != 6'h0);
  assign when_ArraySlice_l113_228 = (7'h40 <= _zz_when_ArraySlice_l113_228);
  always @(*) begin
    if(when_ArraySlice_l112_228) begin
      if(when_ArraySlice_l113_228) begin
        _zz_when_ArraySlice_l173_228 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_228 = (_zz__zz_when_ArraySlice_l173_228 - _zz__zz_when_ArraySlice_l173_228_3);
      end
    end else begin
      if(when_ArraySlice_l118_228) begin
        _zz_when_ArraySlice_l173_228 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_228 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_228 = (_zz_when_ArraySlice_l118_228 <= wReg);
  assign when_ArraySlice_l173_228 = (_zz_when_ArraySlice_l173_228_1 <= _zz_when_ArraySlice_l173_228_3);
  assign when_ArraySlice_l165_229 = (_zz_when_ArraySlice_l165_229 <= selectWriteFifo);
  assign when_ArraySlice_l166_229 = (_zz_when_ArraySlice_l166_229 <= _zz_when_ArraySlice_l166_229_2);
  assign _zz_when_ArraySlice_l112_229 = (wReg % _zz__zz_when_ArraySlice_l112_229);
  assign when_ArraySlice_l112_229 = (_zz_when_ArraySlice_l112_229 != 6'h0);
  assign when_ArraySlice_l113_229 = (7'h40 <= _zz_when_ArraySlice_l113_229);
  always @(*) begin
    if(when_ArraySlice_l112_229) begin
      if(when_ArraySlice_l113_229) begin
        _zz_when_ArraySlice_l173_229 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_229 = (_zz__zz_when_ArraySlice_l173_229 - _zz__zz_when_ArraySlice_l173_229_3);
      end
    end else begin
      if(when_ArraySlice_l118_229) begin
        _zz_when_ArraySlice_l173_229 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_229 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_229 = (_zz_when_ArraySlice_l118_229 <= wReg);
  assign when_ArraySlice_l173_229 = (_zz_when_ArraySlice_l173_229_1 <= _zz_when_ArraySlice_l173_229_3);
  assign when_ArraySlice_l165_230 = (_zz_when_ArraySlice_l165_230 <= selectWriteFifo);
  assign when_ArraySlice_l166_230 = (_zz_when_ArraySlice_l166_230 <= _zz_when_ArraySlice_l166_230_2);
  assign _zz_when_ArraySlice_l112_230 = (wReg % _zz__zz_when_ArraySlice_l112_230);
  assign when_ArraySlice_l112_230 = (_zz_when_ArraySlice_l112_230 != 6'h0);
  assign when_ArraySlice_l113_230 = (7'h40 <= _zz_when_ArraySlice_l113_230);
  always @(*) begin
    if(when_ArraySlice_l112_230) begin
      if(when_ArraySlice_l113_230) begin
        _zz_when_ArraySlice_l173_230 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_230 = (_zz__zz_when_ArraySlice_l173_230 - _zz__zz_when_ArraySlice_l173_230_3);
      end
    end else begin
      if(when_ArraySlice_l118_230) begin
        _zz_when_ArraySlice_l173_230 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_230 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_230 = (_zz_when_ArraySlice_l118_230 <= wReg);
  assign when_ArraySlice_l173_230 = (_zz_when_ArraySlice_l173_230_1 <= _zz_when_ArraySlice_l173_230_3);
  assign when_ArraySlice_l165_231 = (_zz_when_ArraySlice_l165_231 <= selectWriteFifo);
  assign when_ArraySlice_l166_231 = (_zz_when_ArraySlice_l166_231 <= _zz_when_ArraySlice_l166_231_2);
  assign _zz_when_ArraySlice_l112_231 = (wReg % _zz__zz_when_ArraySlice_l112_231);
  assign when_ArraySlice_l112_231 = (_zz_when_ArraySlice_l112_231 != 6'h0);
  assign when_ArraySlice_l113_231 = (7'h40 <= _zz_when_ArraySlice_l113_231);
  always @(*) begin
    if(when_ArraySlice_l112_231) begin
      if(when_ArraySlice_l113_231) begin
        _zz_when_ArraySlice_l173_231 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_231 = (_zz__zz_when_ArraySlice_l173_231 - _zz__zz_when_ArraySlice_l173_231_3);
      end
    end else begin
      if(when_ArraySlice_l118_231) begin
        _zz_when_ArraySlice_l173_231 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_231 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_231 = (_zz_when_ArraySlice_l118_231 <= wReg);
  assign when_ArraySlice_l173_231 = (_zz_when_ArraySlice_l173_231_1 <= _zz_when_ArraySlice_l173_231_3);
  assign when_ArraySlice_l311 = (! ((((((_zz_when_ArraySlice_l311 && _zz_when_ArraySlice_l311_1) && (holdReadOp_4 == _zz_when_ArraySlice_l311_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l311_3 && _zz_when_ArraySlice_l311_4) && (debug_4_28 == _zz_when_ArraySlice_l311_5)) && (debug_5_28 == 1'b1)) && (debug_6_28 == 1'b1)) && (debug_7_28 == 1'b1))));
  assign outputStreamArrayData_0_fire_12 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l315 = ((_zz_when_ArraySlice_l315 == 13'h0) && outputStreamArrayData_0_fire_12);
  assign when_ArraySlice_l301 = (allowPadding_0 && (wReg <= _zz_when_ArraySlice_l301));
  assign outputStreamArrayData_0_fire_13 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l322 = (handshakeTimes_0_value == _zz_when_ArraySlice_l322);
  assign when_ArraySlice_l240_1 = (_zz_when_ArraySlice_l240_1_1 < wReg);
  assign when_ArraySlice_l241_1 = ((! holdReadOp_1) && (_zz_when_ArraySlice_l241_1_1 != 7'h0));
  assign _zz_outputStreamArrayData_1_valid_1 = (selectReadFifo_1 + _zz__zz_outputStreamArrayData_1_valid_1_1);
  assign _zz_12 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_1_valid_1);
  assign _zz_io_pop_ready_9 = outputStreamArrayData_1_ready;
  assign when_ArraySlice_l246_1 = (! holdReadOp_1);
  assign outputStreamArrayData_1_fire_7 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l247_1 = ((_zz_when_ArraySlice_l247_1_1 < _zz_when_ArraySlice_l247_1_3) && outputStreamArrayData_1_fire_7);
  assign when_ArraySlice_l248_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l248_1_1);
  assign when_ArraySlice_l251_1 = (_zz_when_ArraySlice_l251_1_1 == 13'h0);
  assign outputStreamArrayData_1_fire_8 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l256_1 = ((_zz_when_ArraySlice_l256_1_1 == _zz_when_ArraySlice_l256_1_5) && outputStreamArrayData_1_fire_8);
  assign when_ArraySlice_l257_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l257_1_1);
  assign _zz_when_ArraySlice_l94_27 = (hReg % _zz__zz_when_ArraySlice_l94_27);
  assign when_ArraySlice_l94_27 = (_zz_when_ArraySlice_l94_27 != 6'h0);
  assign when_ArraySlice_l95_27 = (7'h40 <= _zz_when_ArraySlice_l95_27);
  always @(*) begin
    if(when_ArraySlice_l94_27) begin
      if(when_ArraySlice_l95_27) begin
        _zz_when_ArraySlice_l259_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_1 = (_zz__zz_when_ArraySlice_l259_1_1 - _zz__zz_when_ArraySlice_l259_1_4);
      end
    end else begin
      if(when_ArraySlice_l99_27) begin
        _zz_when_ArraySlice_l259_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_1 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_27 = (_zz_when_ArraySlice_l99_27 <= hReg);
  assign when_ArraySlice_l259_1 = (_zz_when_ArraySlice_l259_1_1 < _zz_when_ArraySlice_l259_1_4);
  always @(*) begin
    debug_0_29 = 1'b0;
    if(when_ArraySlice_l165_232) begin
      if(when_ArraySlice_l166_232) begin
        debug_0_29 = 1'b1;
      end else begin
        debug_0_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_232) begin
        debug_0_29 = 1'b1;
      end else begin
        debug_0_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_29 = 1'b0;
    if(when_ArraySlice_l165_233) begin
      if(when_ArraySlice_l166_233) begin
        debug_1_29 = 1'b1;
      end else begin
        debug_1_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_233) begin
        debug_1_29 = 1'b1;
      end else begin
        debug_1_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_29 = 1'b0;
    if(when_ArraySlice_l165_234) begin
      if(when_ArraySlice_l166_234) begin
        debug_2_29 = 1'b1;
      end else begin
        debug_2_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_234) begin
        debug_2_29 = 1'b1;
      end else begin
        debug_2_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_29 = 1'b0;
    if(when_ArraySlice_l165_235) begin
      if(when_ArraySlice_l166_235) begin
        debug_3_29 = 1'b1;
      end else begin
        debug_3_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_235) begin
        debug_3_29 = 1'b1;
      end else begin
        debug_3_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_29 = 1'b0;
    if(when_ArraySlice_l165_236) begin
      if(when_ArraySlice_l166_236) begin
        debug_4_29 = 1'b1;
      end else begin
        debug_4_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_236) begin
        debug_4_29 = 1'b1;
      end else begin
        debug_4_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_29 = 1'b0;
    if(when_ArraySlice_l165_237) begin
      if(when_ArraySlice_l166_237) begin
        debug_5_29 = 1'b1;
      end else begin
        debug_5_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_237) begin
        debug_5_29 = 1'b1;
      end else begin
        debug_5_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_29 = 1'b0;
    if(when_ArraySlice_l165_238) begin
      if(when_ArraySlice_l166_238) begin
        debug_6_29 = 1'b1;
      end else begin
        debug_6_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_238) begin
        debug_6_29 = 1'b1;
      end else begin
        debug_6_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_29 = 1'b0;
    if(when_ArraySlice_l165_239) begin
      if(when_ArraySlice_l166_239) begin
        debug_7_29 = 1'b1;
      end else begin
        debug_7_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_239) begin
        debug_7_29 = 1'b1;
      end else begin
        debug_7_29 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_232 = (_zz_when_ArraySlice_l165_232 <= selectWriteFifo);
  assign when_ArraySlice_l166_232 = (_zz_when_ArraySlice_l166_232 <= _zz_when_ArraySlice_l166_232_1);
  assign _zz_when_ArraySlice_l112_232 = (wReg % _zz__zz_when_ArraySlice_l112_232);
  assign when_ArraySlice_l112_232 = (_zz_when_ArraySlice_l112_232 != 6'h0);
  assign when_ArraySlice_l113_232 = (7'h40 <= _zz_when_ArraySlice_l113_232);
  always @(*) begin
    if(when_ArraySlice_l112_232) begin
      if(when_ArraySlice_l113_232) begin
        _zz_when_ArraySlice_l173_232 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_232 = (_zz__zz_when_ArraySlice_l173_232 - _zz__zz_when_ArraySlice_l173_232_3);
      end
    end else begin
      if(when_ArraySlice_l118_232) begin
        _zz_when_ArraySlice_l173_232 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_232 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_232 = (_zz_when_ArraySlice_l118_232 <= wReg);
  assign when_ArraySlice_l173_232 = (_zz_when_ArraySlice_l173_232_1 <= _zz_when_ArraySlice_l173_232_2);
  assign when_ArraySlice_l165_233 = (_zz_when_ArraySlice_l165_233 <= selectWriteFifo);
  assign when_ArraySlice_l166_233 = (_zz_when_ArraySlice_l166_233 <= _zz_when_ArraySlice_l166_233_1);
  assign _zz_when_ArraySlice_l112_233 = (wReg % _zz__zz_when_ArraySlice_l112_233);
  assign when_ArraySlice_l112_233 = (_zz_when_ArraySlice_l112_233 != 6'h0);
  assign when_ArraySlice_l113_233 = (7'h40 <= _zz_when_ArraySlice_l113_233);
  always @(*) begin
    if(when_ArraySlice_l112_233) begin
      if(when_ArraySlice_l113_233) begin
        _zz_when_ArraySlice_l173_233 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_233 = (_zz__zz_when_ArraySlice_l173_233 - _zz__zz_when_ArraySlice_l173_233_3);
      end
    end else begin
      if(when_ArraySlice_l118_233) begin
        _zz_when_ArraySlice_l173_233 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_233 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_233 = (_zz_when_ArraySlice_l118_233 <= wReg);
  assign when_ArraySlice_l173_233 = (_zz_when_ArraySlice_l173_233_1 <= _zz_when_ArraySlice_l173_233_3);
  assign when_ArraySlice_l165_234 = (_zz_when_ArraySlice_l165_234 <= selectWriteFifo);
  assign when_ArraySlice_l166_234 = (_zz_when_ArraySlice_l166_234 <= _zz_when_ArraySlice_l166_234_1);
  assign _zz_when_ArraySlice_l112_234 = (wReg % _zz__zz_when_ArraySlice_l112_234);
  assign when_ArraySlice_l112_234 = (_zz_when_ArraySlice_l112_234 != 6'h0);
  assign when_ArraySlice_l113_234 = (7'h40 <= _zz_when_ArraySlice_l113_234);
  always @(*) begin
    if(when_ArraySlice_l112_234) begin
      if(when_ArraySlice_l113_234) begin
        _zz_when_ArraySlice_l173_234 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_234 = (_zz__zz_when_ArraySlice_l173_234 - _zz__zz_when_ArraySlice_l173_234_3);
      end
    end else begin
      if(when_ArraySlice_l118_234) begin
        _zz_when_ArraySlice_l173_234 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_234 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_234 = (_zz_when_ArraySlice_l118_234 <= wReg);
  assign when_ArraySlice_l173_234 = (_zz_when_ArraySlice_l173_234_1 <= _zz_when_ArraySlice_l173_234_3);
  assign when_ArraySlice_l165_235 = (_zz_when_ArraySlice_l165_235 <= selectWriteFifo);
  assign when_ArraySlice_l166_235 = (_zz_when_ArraySlice_l166_235 <= _zz_when_ArraySlice_l166_235_1);
  assign _zz_when_ArraySlice_l112_235 = (wReg % _zz__zz_when_ArraySlice_l112_235);
  assign when_ArraySlice_l112_235 = (_zz_when_ArraySlice_l112_235 != 6'h0);
  assign when_ArraySlice_l113_235 = (7'h40 <= _zz_when_ArraySlice_l113_235);
  always @(*) begin
    if(when_ArraySlice_l112_235) begin
      if(when_ArraySlice_l113_235) begin
        _zz_when_ArraySlice_l173_235 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_235 = (_zz__zz_when_ArraySlice_l173_235 - _zz__zz_when_ArraySlice_l173_235_3);
      end
    end else begin
      if(when_ArraySlice_l118_235) begin
        _zz_when_ArraySlice_l173_235 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_235 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_235 = (_zz_when_ArraySlice_l118_235 <= wReg);
  assign when_ArraySlice_l173_235 = (_zz_when_ArraySlice_l173_235_1 <= _zz_when_ArraySlice_l173_235_3);
  assign when_ArraySlice_l165_236 = (_zz_when_ArraySlice_l165_236 <= selectWriteFifo);
  assign when_ArraySlice_l166_236 = (_zz_when_ArraySlice_l166_236 <= _zz_when_ArraySlice_l166_236_1);
  assign _zz_when_ArraySlice_l112_236 = (wReg % _zz__zz_when_ArraySlice_l112_236);
  assign when_ArraySlice_l112_236 = (_zz_when_ArraySlice_l112_236 != 6'h0);
  assign when_ArraySlice_l113_236 = (7'h40 <= _zz_when_ArraySlice_l113_236);
  always @(*) begin
    if(when_ArraySlice_l112_236) begin
      if(when_ArraySlice_l113_236) begin
        _zz_when_ArraySlice_l173_236 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_236 = (_zz__zz_when_ArraySlice_l173_236 - _zz__zz_when_ArraySlice_l173_236_3);
      end
    end else begin
      if(when_ArraySlice_l118_236) begin
        _zz_when_ArraySlice_l173_236 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_236 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_236 = (_zz_when_ArraySlice_l118_236 <= wReg);
  assign when_ArraySlice_l173_236 = (_zz_when_ArraySlice_l173_236_1 <= _zz_when_ArraySlice_l173_236_3);
  assign when_ArraySlice_l165_237 = (_zz_when_ArraySlice_l165_237 <= selectWriteFifo);
  assign when_ArraySlice_l166_237 = (_zz_when_ArraySlice_l166_237 <= _zz_when_ArraySlice_l166_237_2);
  assign _zz_when_ArraySlice_l112_237 = (wReg % _zz__zz_when_ArraySlice_l112_237);
  assign when_ArraySlice_l112_237 = (_zz_when_ArraySlice_l112_237 != 6'h0);
  assign when_ArraySlice_l113_237 = (7'h40 <= _zz_when_ArraySlice_l113_237);
  always @(*) begin
    if(when_ArraySlice_l112_237) begin
      if(when_ArraySlice_l113_237) begin
        _zz_when_ArraySlice_l173_237 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_237 = (_zz__zz_when_ArraySlice_l173_237 - _zz__zz_when_ArraySlice_l173_237_3);
      end
    end else begin
      if(when_ArraySlice_l118_237) begin
        _zz_when_ArraySlice_l173_237 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_237 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_237 = (_zz_when_ArraySlice_l118_237 <= wReg);
  assign when_ArraySlice_l173_237 = (_zz_when_ArraySlice_l173_237_1 <= _zz_when_ArraySlice_l173_237_3);
  assign when_ArraySlice_l165_238 = (_zz_when_ArraySlice_l165_238 <= selectWriteFifo);
  assign when_ArraySlice_l166_238 = (_zz_when_ArraySlice_l166_238 <= _zz_when_ArraySlice_l166_238_2);
  assign _zz_when_ArraySlice_l112_238 = (wReg % _zz__zz_when_ArraySlice_l112_238);
  assign when_ArraySlice_l112_238 = (_zz_when_ArraySlice_l112_238 != 6'h0);
  assign when_ArraySlice_l113_238 = (7'h40 <= _zz_when_ArraySlice_l113_238);
  always @(*) begin
    if(when_ArraySlice_l112_238) begin
      if(when_ArraySlice_l113_238) begin
        _zz_when_ArraySlice_l173_238 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_238 = (_zz__zz_when_ArraySlice_l173_238 - _zz__zz_when_ArraySlice_l173_238_3);
      end
    end else begin
      if(when_ArraySlice_l118_238) begin
        _zz_when_ArraySlice_l173_238 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_238 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_238 = (_zz_when_ArraySlice_l118_238 <= wReg);
  assign when_ArraySlice_l173_238 = (_zz_when_ArraySlice_l173_238_1 <= _zz_when_ArraySlice_l173_238_3);
  assign when_ArraySlice_l165_239 = (_zz_when_ArraySlice_l165_239 <= selectWriteFifo);
  assign when_ArraySlice_l166_239 = (_zz_when_ArraySlice_l166_239 <= _zz_when_ArraySlice_l166_239_2);
  assign _zz_when_ArraySlice_l112_239 = (wReg % _zz__zz_when_ArraySlice_l112_239);
  assign when_ArraySlice_l112_239 = (_zz_when_ArraySlice_l112_239 != 6'h0);
  assign when_ArraySlice_l113_239 = (7'h40 <= _zz_when_ArraySlice_l113_239);
  always @(*) begin
    if(when_ArraySlice_l112_239) begin
      if(when_ArraySlice_l113_239) begin
        _zz_when_ArraySlice_l173_239 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_239 = (_zz__zz_when_ArraySlice_l173_239 - _zz__zz_when_ArraySlice_l173_239_3);
      end
    end else begin
      if(when_ArraySlice_l118_239) begin
        _zz_when_ArraySlice_l173_239 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_239 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_239 = (_zz_when_ArraySlice_l118_239 <= wReg);
  assign when_ArraySlice_l173_239 = (_zz_when_ArraySlice_l173_239_1 <= _zz_when_ArraySlice_l173_239_3);
  assign when_ArraySlice_l265_1 = (! ((((((_zz_when_ArraySlice_l265_1_1 && _zz_when_ArraySlice_l265_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l265_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l265_1_4 && _zz_when_ArraySlice_l265_1_5) && (debug_4_29 == _zz_when_ArraySlice_l265_1_6)) && (debug_5_29 == 1'b1)) && (debug_6_29 == 1'b1)) && (debug_7_29 == 1'b1))));
  assign when_ArraySlice_l268_1 = (wReg <= _zz_when_ArraySlice_l268_1_1);
  assign when_ArraySlice_l272_1 = (_zz_when_ArraySlice_l272_1_1 == 13'h0);
  assign when_ArraySlice_l276_1 = (_zz_when_ArraySlice_l276_1_1 == 7'h0);
  assign outputStreamArrayData_1_fire_9 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l277_1 = ((handshakeTimes_1_value == _zz_when_ArraySlice_l277_1_1) && outputStreamArrayData_1_fire_9);
  assign _zz_when_ArraySlice_l94_28 = (hReg % _zz__zz_when_ArraySlice_l94_28);
  assign when_ArraySlice_l94_28 = (_zz_when_ArraySlice_l94_28 != 6'h0);
  assign when_ArraySlice_l95_28 = (7'h40 <= _zz_when_ArraySlice_l95_28);
  always @(*) begin
    if(when_ArraySlice_l94_28) begin
      if(when_ArraySlice_l95_28) begin
        _zz_when_ArraySlice_l279_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_1 = (_zz__zz_when_ArraySlice_l279_1_1 - _zz__zz_when_ArraySlice_l279_1_4);
      end
    end else begin
      if(when_ArraySlice_l99_28) begin
        _zz_when_ArraySlice_l279_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_1 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_28 = (_zz_when_ArraySlice_l99_28 <= hReg);
  assign when_ArraySlice_l279_1 = (_zz_when_ArraySlice_l279_1_1 < _zz_when_ArraySlice_l279_1_4);
  always @(*) begin
    debug_0_30 = 1'b0;
    if(when_ArraySlice_l165_240) begin
      if(when_ArraySlice_l166_240) begin
        debug_0_30 = 1'b1;
      end else begin
        debug_0_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_240) begin
        debug_0_30 = 1'b1;
      end else begin
        debug_0_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_30 = 1'b0;
    if(when_ArraySlice_l165_241) begin
      if(when_ArraySlice_l166_241) begin
        debug_1_30 = 1'b1;
      end else begin
        debug_1_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_241) begin
        debug_1_30 = 1'b1;
      end else begin
        debug_1_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_30 = 1'b0;
    if(when_ArraySlice_l165_242) begin
      if(when_ArraySlice_l166_242) begin
        debug_2_30 = 1'b1;
      end else begin
        debug_2_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_242) begin
        debug_2_30 = 1'b1;
      end else begin
        debug_2_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_30 = 1'b0;
    if(when_ArraySlice_l165_243) begin
      if(when_ArraySlice_l166_243) begin
        debug_3_30 = 1'b1;
      end else begin
        debug_3_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_243) begin
        debug_3_30 = 1'b1;
      end else begin
        debug_3_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_30 = 1'b0;
    if(when_ArraySlice_l165_244) begin
      if(when_ArraySlice_l166_244) begin
        debug_4_30 = 1'b1;
      end else begin
        debug_4_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_244) begin
        debug_4_30 = 1'b1;
      end else begin
        debug_4_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_30 = 1'b0;
    if(when_ArraySlice_l165_245) begin
      if(when_ArraySlice_l166_245) begin
        debug_5_30 = 1'b1;
      end else begin
        debug_5_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_245) begin
        debug_5_30 = 1'b1;
      end else begin
        debug_5_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_30 = 1'b0;
    if(when_ArraySlice_l165_246) begin
      if(when_ArraySlice_l166_246) begin
        debug_6_30 = 1'b1;
      end else begin
        debug_6_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_246) begin
        debug_6_30 = 1'b1;
      end else begin
        debug_6_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_30 = 1'b0;
    if(when_ArraySlice_l165_247) begin
      if(when_ArraySlice_l166_247) begin
        debug_7_30 = 1'b1;
      end else begin
        debug_7_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_247) begin
        debug_7_30 = 1'b1;
      end else begin
        debug_7_30 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_240 = (_zz_when_ArraySlice_l165_240 <= selectWriteFifo);
  assign when_ArraySlice_l166_240 = (_zz_when_ArraySlice_l166_240 <= _zz_when_ArraySlice_l166_240_1);
  assign _zz_when_ArraySlice_l112_240 = (wReg % _zz__zz_when_ArraySlice_l112_240);
  assign when_ArraySlice_l112_240 = (_zz_when_ArraySlice_l112_240 != 6'h0);
  assign when_ArraySlice_l113_240 = (7'h40 <= _zz_when_ArraySlice_l113_240);
  always @(*) begin
    if(when_ArraySlice_l112_240) begin
      if(when_ArraySlice_l113_240) begin
        _zz_when_ArraySlice_l173_240 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_240 = (_zz__zz_when_ArraySlice_l173_240 - _zz__zz_when_ArraySlice_l173_240_3);
      end
    end else begin
      if(when_ArraySlice_l118_240) begin
        _zz_when_ArraySlice_l173_240 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_240 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_240 = (_zz_when_ArraySlice_l118_240 <= wReg);
  assign when_ArraySlice_l173_240 = (_zz_when_ArraySlice_l173_240_1 <= _zz_when_ArraySlice_l173_240_2);
  assign when_ArraySlice_l165_241 = (_zz_when_ArraySlice_l165_241 <= selectWriteFifo);
  assign when_ArraySlice_l166_241 = (_zz_when_ArraySlice_l166_241 <= _zz_when_ArraySlice_l166_241_1);
  assign _zz_when_ArraySlice_l112_241 = (wReg % _zz__zz_when_ArraySlice_l112_241);
  assign when_ArraySlice_l112_241 = (_zz_when_ArraySlice_l112_241 != 6'h0);
  assign when_ArraySlice_l113_241 = (7'h40 <= _zz_when_ArraySlice_l113_241);
  always @(*) begin
    if(when_ArraySlice_l112_241) begin
      if(when_ArraySlice_l113_241) begin
        _zz_when_ArraySlice_l173_241 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_241 = (_zz__zz_when_ArraySlice_l173_241 - _zz__zz_when_ArraySlice_l173_241_3);
      end
    end else begin
      if(when_ArraySlice_l118_241) begin
        _zz_when_ArraySlice_l173_241 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_241 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_241 = (_zz_when_ArraySlice_l118_241 <= wReg);
  assign when_ArraySlice_l173_241 = (_zz_when_ArraySlice_l173_241_1 <= _zz_when_ArraySlice_l173_241_3);
  assign when_ArraySlice_l165_242 = (_zz_when_ArraySlice_l165_242 <= selectWriteFifo);
  assign when_ArraySlice_l166_242 = (_zz_when_ArraySlice_l166_242 <= _zz_when_ArraySlice_l166_242_1);
  assign _zz_when_ArraySlice_l112_242 = (wReg % _zz__zz_when_ArraySlice_l112_242);
  assign when_ArraySlice_l112_242 = (_zz_when_ArraySlice_l112_242 != 6'h0);
  assign when_ArraySlice_l113_242 = (7'h40 <= _zz_when_ArraySlice_l113_242);
  always @(*) begin
    if(when_ArraySlice_l112_242) begin
      if(when_ArraySlice_l113_242) begin
        _zz_when_ArraySlice_l173_242 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_242 = (_zz__zz_when_ArraySlice_l173_242 - _zz__zz_when_ArraySlice_l173_242_3);
      end
    end else begin
      if(when_ArraySlice_l118_242) begin
        _zz_when_ArraySlice_l173_242 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_242 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_242 = (_zz_when_ArraySlice_l118_242 <= wReg);
  assign when_ArraySlice_l173_242 = (_zz_when_ArraySlice_l173_242_1 <= _zz_when_ArraySlice_l173_242_3);
  assign when_ArraySlice_l165_243 = (_zz_when_ArraySlice_l165_243 <= selectWriteFifo);
  assign when_ArraySlice_l166_243 = (_zz_when_ArraySlice_l166_243 <= _zz_when_ArraySlice_l166_243_1);
  assign _zz_when_ArraySlice_l112_243 = (wReg % _zz__zz_when_ArraySlice_l112_243);
  assign when_ArraySlice_l112_243 = (_zz_when_ArraySlice_l112_243 != 6'h0);
  assign when_ArraySlice_l113_243 = (7'h40 <= _zz_when_ArraySlice_l113_243);
  always @(*) begin
    if(when_ArraySlice_l112_243) begin
      if(when_ArraySlice_l113_243) begin
        _zz_when_ArraySlice_l173_243 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_243 = (_zz__zz_when_ArraySlice_l173_243 - _zz__zz_when_ArraySlice_l173_243_3);
      end
    end else begin
      if(when_ArraySlice_l118_243) begin
        _zz_when_ArraySlice_l173_243 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_243 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_243 = (_zz_when_ArraySlice_l118_243 <= wReg);
  assign when_ArraySlice_l173_243 = (_zz_when_ArraySlice_l173_243_1 <= _zz_when_ArraySlice_l173_243_3);
  assign when_ArraySlice_l165_244 = (_zz_when_ArraySlice_l165_244 <= selectWriteFifo);
  assign when_ArraySlice_l166_244 = (_zz_when_ArraySlice_l166_244 <= _zz_when_ArraySlice_l166_244_1);
  assign _zz_when_ArraySlice_l112_244 = (wReg % _zz__zz_when_ArraySlice_l112_244);
  assign when_ArraySlice_l112_244 = (_zz_when_ArraySlice_l112_244 != 6'h0);
  assign when_ArraySlice_l113_244 = (7'h40 <= _zz_when_ArraySlice_l113_244);
  always @(*) begin
    if(when_ArraySlice_l112_244) begin
      if(when_ArraySlice_l113_244) begin
        _zz_when_ArraySlice_l173_244 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_244 = (_zz__zz_when_ArraySlice_l173_244 - _zz__zz_when_ArraySlice_l173_244_3);
      end
    end else begin
      if(when_ArraySlice_l118_244) begin
        _zz_when_ArraySlice_l173_244 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_244 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_244 = (_zz_when_ArraySlice_l118_244 <= wReg);
  assign when_ArraySlice_l173_244 = (_zz_when_ArraySlice_l173_244_1 <= _zz_when_ArraySlice_l173_244_3);
  assign when_ArraySlice_l165_245 = (_zz_when_ArraySlice_l165_245 <= selectWriteFifo);
  assign when_ArraySlice_l166_245 = (_zz_when_ArraySlice_l166_245 <= _zz_when_ArraySlice_l166_245_2);
  assign _zz_when_ArraySlice_l112_245 = (wReg % _zz__zz_when_ArraySlice_l112_245);
  assign when_ArraySlice_l112_245 = (_zz_when_ArraySlice_l112_245 != 6'h0);
  assign when_ArraySlice_l113_245 = (7'h40 <= _zz_when_ArraySlice_l113_245);
  always @(*) begin
    if(when_ArraySlice_l112_245) begin
      if(when_ArraySlice_l113_245) begin
        _zz_when_ArraySlice_l173_245 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_245 = (_zz__zz_when_ArraySlice_l173_245 - _zz__zz_when_ArraySlice_l173_245_3);
      end
    end else begin
      if(when_ArraySlice_l118_245) begin
        _zz_when_ArraySlice_l173_245 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_245 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_245 = (_zz_when_ArraySlice_l118_245 <= wReg);
  assign when_ArraySlice_l173_245 = (_zz_when_ArraySlice_l173_245_1 <= _zz_when_ArraySlice_l173_245_3);
  assign when_ArraySlice_l165_246 = (_zz_when_ArraySlice_l165_246 <= selectWriteFifo);
  assign when_ArraySlice_l166_246 = (_zz_when_ArraySlice_l166_246 <= _zz_when_ArraySlice_l166_246_2);
  assign _zz_when_ArraySlice_l112_246 = (wReg % _zz__zz_when_ArraySlice_l112_246);
  assign when_ArraySlice_l112_246 = (_zz_when_ArraySlice_l112_246 != 6'h0);
  assign when_ArraySlice_l113_246 = (7'h40 <= _zz_when_ArraySlice_l113_246);
  always @(*) begin
    if(when_ArraySlice_l112_246) begin
      if(when_ArraySlice_l113_246) begin
        _zz_when_ArraySlice_l173_246 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_246 = (_zz__zz_when_ArraySlice_l173_246 - _zz__zz_when_ArraySlice_l173_246_3);
      end
    end else begin
      if(when_ArraySlice_l118_246) begin
        _zz_when_ArraySlice_l173_246 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_246 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_246 = (_zz_when_ArraySlice_l118_246 <= wReg);
  assign when_ArraySlice_l173_246 = (_zz_when_ArraySlice_l173_246_1 <= _zz_when_ArraySlice_l173_246_3);
  assign when_ArraySlice_l165_247 = (_zz_when_ArraySlice_l165_247 <= selectWriteFifo);
  assign when_ArraySlice_l166_247 = (_zz_when_ArraySlice_l166_247 <= _zz_when_ArraySlice_l166_247_2);
  assign _zz_when_ArraySlice_l112_247 = (wReg % _zz__zz_when_ArraySlice_l112_247);
  assign when_ArraySlice_l112_247 = (_zz_when_ArraySlice_l112_247 != 6'h0);
  assign when_ArraySlice_l113_247 = (7'h40 <= _zz_when_ArraySlice_l113_247);
  always @(*) begin
    if(when_ArraySlice_l112_247) begin
      if(when_ArraySlice_l113_247) begin
        _zz_when_ArraySlice_l173_247 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_247 = (_zz__zz_when_ArraySlice_l173_247 - _zz__zz_when_ArraySlice_l173_247_3);
      end
    end else begin
      if(when_ArraySlice_l118_247) begin
        _zz_when_ArraySlice_l173_247 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_247 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_247 = (_zz_when_ArraySlice_l118_247 <= wReg);
  assign when_ArraySlice_l173_247 = (_zz_when_ArraySlice_l173_247_1 <= _zz_when_ArraySlice_l173_247_3);
  assign when_ArraySlice_l285_1 = (! ((((((_zz_when_ArraySlice_l285_1_1 && _zz_when_ArraySlice_l285_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l285_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l285_1_4 && _zz_when_ArraySlice_l285_1_5) && (debug_4_30 == _zz_when_ArraySlice_l285_1_6)) && (debug_5_30 == 1'b1)) && (debug_6_30 == 1'b1)) && (debug_7_30 == 1'b1))));
  assign when_ArraySlice_l288_1 = (wReg <= _zz_when_ArraySlice_l288_1_1);
  assign outputStreamArrayData_1_fire_10 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l292_1 = ((_zz_when_ArraySlice_l292_1_1 == 13'h0) && outputStreamArrayData_1_fire_10);
  assign outputStreamArrayData_1_fire_11 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l303_1 = ((handshakeTimes_1_value == _zz_when_ArraySlice_l303_1_1) && outputStreamArrayData_1_fire_11);
  assign _zz_when_ArraySlice_l94_29 = (hReg % _zz__zz_when_ArraySlice_l94_29);
  assign when_ArraySlice_l94_29 = (_zz_when_ArraySlice_l94_29 != 6'h0);
  assign when_ArraySlice_l95_29 = (7'h40 <= _zz_when_ArraySlice_l95_29);
  always @(*) begin
    if(when_ArraySlice_l94_29) begin
      if(when_ArraySlice_l95_29) begin
        _zz_when_ArraySlice_l304_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_1 = (_zz__zz_when_ArraySlice_l304_1_1 - _zz__zz_when_ArraySlice_l304_1_4);
      end
    end else begin
      if(when_ArraySlice_l99_29) begin
        _zz_when_ArraySlice_l304_1 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_1 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_29 = (_zz_when_ArraySlice_l99_29 <= hReg);
  assign when_ArraySlice_l304_1 = (_zz_when_ArraySlice_l304_1_1 < _zz_when_ArraySlice_l304_1_4);
  always @(*) begin
    debug_0_31 = 1'b0;
    if(when_ArraySlice_l165_248) begin
      if(when_ArraySlice_l166_248) begin
        debug_0_31 = 1'b1;
      end else begin
        debug_0_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_248) begin
        debug_0_31 = 1'b1;
      end else begin
        debug_0_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_31 = 1'b0;
    if(when_ArraySlice_l165_249) begin
      if(when_ArraySlice_l166_249) begin
        debug_1_31 = 1'b1;
      end else begin
        debug_1_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_249) begin
        debug_1_31 = 1'b1;
      end else begin
        debug_1_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_31 = 1'b0;
    if(when_ArraySlice_l165_250) begin
      if(when_ArraySlice_l166_250) begin
        debug_2_31 = 1'b1;
      end else begin
        debug_2_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_250) begin
        debug_2_31 = 1'b1;
      end else begin
        debug_2_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_31 = 1'b0;
    if(when_ArraySlice_l165_251) begin
      if(when_ArraySlice_l166_251) begin
        debug_3_31 = 1'b1;
      end else begin
        debug_3_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_251) begin
        debug_3_31 = 1'b1;
      end else begin
        debug_3_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_31 = 1'b0;
    if(when_ArraySlice_l165_252) begin
      if(when_ArraySlice_l166_252) begin
        debug_4_31 = 1'b1;
      end else begin
        debug_4_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_252) begin
        debug_4_31 = 1'b1;
      end else begin
        debug_4_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_31 = 1'b0;
    if(when_ArraySlice_l165_253) begin
      if(when_ArraySlice_l166_253) begin
        debug_5_31 = 1'b1;
      end else begin
        debug_5_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_253) begin
        debug_5_31 = 1'b1;
      end else begin
        debug_5_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_31 = 1'b0;
    if(when_ArraySlice_l165_254) begin
      if(when_ArraySlice_l166_254) begin
        debug_6_31 = 1'b1;
      end else begin
        debug_6_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_254) begin
        debug_6_31 = 1'b1;
      end else begin
        debug_6_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_31 = 1'b0;
    if(when_ArraySlice_l165_255) begin
      if(when_ArraySlice_l166_255) begin
        debug_7_31 = 1'b1;
      end else begin
        debug_7_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_255) begin
        debug_7_31 = 1'b1;
      end else begin
        debug_7_31 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_248 = (_zz_when_ArraySlice_l165_248 <= selectWriteFifo);
  assign when_ArraySlice_l166_248 = (_zz_when_ArraySlice_l166_248 <= _zz_when_ArraySlice_l166_248_1);
  assign _zz_when_ArraySlice_l112_248 = (wReg % _zz__zz_when_ArraySlice_l112_248);
  assign when_ArraySlice_l112_248 = (_zz_when_ArraySlice_l112_248 != 6'h0);
  assign when_ArraySlice_l113_248 = (7'h40 <= _zz_when_ArraySlice_l113_248);
  always @(*) begin
    if(when_ArraySlice_l112_248) begin
      if(when_ArraySlice_l113_248) begin
        _zz_when_ArraySlice_l173_248 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_248 = (_zz__zz_when_ArraySlice_l173_248 - _zz__zz_when_ArraySlice_l173_248_3);
      end
    end else begin
      if(when_ArraySlice_l118_248) begin
        _zz_when_ArraySlice_l173_248 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_248 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_248 = (_zz_when_ArraySlice_l118_248 <= wReg);
  assign when_ArraySlice_l173_248 = (_zz_when_ArraySlice_l173_248_1 <= _zz_when_ArraySlice_l173_248_2);
  assign when_ArraySlice_l165_249 = (_zz_when_ArraySlice_l165_249 <= selectWriteFifo);
  assign when_ArraySlice_l166_249 = (_zz_when_ArraySlice_l166_249 <= _zz_when_ArraySlice_l166_249_1);
  assign _zz_when_ArraySlice_l112_249 = (wReg % _zz__zz_when_ArraySlice_l112_249);
  assign when_ArraySlice_l112_249 = (_zz_when_ArraySlice_l112_249 != 6'h0);
  assign when_ArraySlice_l113_249 = (7'h40 <= _zz_when_ArraySlice_l113_249);
  always @(*) begin
    if(when_ArraySlice_l112_249) begin
      if(when_ArraySlice_l113_249) begin
        _zz_when_ArraySlice_l173_249 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_249 = (_zz__zz_when_ArraySlice_l173_249 - _zz__zz_when_ArraySlice_l173_249_3);
      end
    end else begin
      if(when_ArraySlice_l118_249) begin
        _zz_when_ArraySlice_l173_249 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_249 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_249 = (_zz_when_ArraySlice_l118_249 <= wReg);
  assign when_ArraySlice_l173_249 = (_zz_when_ArraySlice_l173_249_1 <= _zz_when_ArraySlice_l173_249_3);
  assign when_ArraySlice_l165_250 = (_zz_when_ArraySlice_l165_250 <= selectWriteFifo);
  assign when_ArraySlice_l166_250 = (_zz_when_ArraySlice_l166_250 <= _zz_when_ArraySlice_l166_250_1);
  assign _zz_when_ArraySlice_l112_250 = (wReg % _zz__zz_when_ArraySlice_l112_250);
  assign when_ArraySlice_l112_250 = (_zz_when_ArraySlice_l112_250 != 6'h0);
  assign when_ArraySlice_l113_250 = (7'h40 <= _zz_when_ArraySlice_l113_250);
  always @(*) begin
    if(when_ArraySlice_l112_250) begin
      if(when_ArraySlice_l113_250) begin
        _zz_when_ArraySlice_l173_250 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_250 = (_zz__zz_when_ArraySlice_l173_250 - _zz__zz_when_ArraySlice_l173_250_3);
      end
    end else begin
      if(when_ArraySlice_l118_250) begin
        _zz_when_ArraySlice_l173_250 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_250 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_250 = (_zz_when_ArraySlice_l118_250 <= wReg);
  assign when_ArraySlice_l173_250 = (_zz_when_ArraySlice_l173_250_1 <= _zz_when_ArraySlice_l173_250_3);
  assign when_ArraySlice_l165_251 = (_zz_when_ArraySlice_l165_251 <= selectWriteFifo);
  assign when_ArraySlice_l166_251 = (_zz_when_ArraySlice_l166_251 <= _zz_when_ArraySlice_l166_251_1);
  assign _zz_when_ArraySlice_l112_251 = (wReg % _zz__zz_when_ArraySlice_l112_251);
  assign when_ArraySlice_l112_251 = (_zz_when_ArraySlice_l112_251 != 6'h0);
  assign when_ArraySlice_l113_251 = (7'h40 <= _zz_when_ArraySlice_l113_251);
  always @(*) begin
    if(when_ArraySlice_l112_251) begin
      if(when_ArraySlice_l113_251) begin
        _zz_when_ArraySlice_l173_251 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_251 = (_zz__zz_when_ArraySlice_l173_251 - _zz__zz_when_ArraySlice_l173_251_3);
      end
    end else begin
      if(when_ArraySlice_l118_251) begin
        _zz_when_ArraySlice_l173_251 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_251 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_251 = (_zz_when_ArraySlice_l118_251 <= wReg);
  assign when_ArraySlice_l173_251 = (_zz_when_ArraySlice_l173_251_1 <= _zz_when_ArraySlice_l173_251_3);
  assign when_ArraySlice_l165_252 = (_zz_when_ArraySlice_l165_252 <= selectWriteFifo);
  assign when_ArraySlice_l166_252 = (_zz_when_ArraySlice_l166_252 <= _zz_when_ArraySlice_l166_252_1);
  assign _zz_when_ArraySlice_l112_252 = (wReg % _zz__zz_when_ArraySlice_l112_252);
  assign when_ArraySlice_l112_252 = (_zz_when_ArraySlice_l112_252 != 6'h0);
  assign when_ArraySlice_l113_252 = (7'h40 <= _zz_when_ArraySlice_l113_252);
  always @(*) begin
    if(when_ArraySlice_l112_252) begin
      if(when_ArraySlice_l113_252) begin
        _zz_when_ArraySlice_l173_252 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_252 = (_zz__zz_when_ArraySlice_l173_252 - _zz__zz_when_ArraySlice_l173_252_3);
      end
    end else begin
      if(when_ArraySlice_l118_252) begin
        _zz_when_ArraySlice_l173_252 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_252 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_252 = (_zz_when_ArraySlice_l118_252 <= wReg);
  assign when_ArraySlice_l173_252 = (_zz_when_ArraySlice_l173_252_1 <= _zz_when_ArraySlice_l173_252_3);
  assign when_ArraySlice_l165_253 = (_zz_when_ArraySlice_l165_253 <= selectWriteFifo);
  assign when_ArraySlice_l166_253 = (_zz_when_ArraySlice_l166_253 <= _zz_when_ArraySlice_l166_253_2);
  assign _zz_when_ArraySlice_l112_253 = (wReg % _zz__zz_when_ArraySlice_l112_253);
  assign when_ArraySlice_l112_253 = (_zz_when_ArraySlice_l112_253 != 6'h0);
  assign when_ArraySlice_l113_253 = (7'h40 <= _zz_when_ArraySlice_l113_253);
  always @(*) begin
    if(when_ArraySlice_l112_253) begin
      if(when_ArraySlice_l113_253) begin
        _zz_when_ArraySlice_l173_253 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_253 = (_zz__zz_when_ArraySlice_l173_253 - _zz__zz_when_ArraySlice_l173_253_3);
      end
    end else begin
      if(when_ArraySlice_l118_253) begin
        _zz_when_ArraySlice_l173_253 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_253 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_253 = (_zz_when_ArraySlice_l118_253 <= wReg);
  assign when_ArraySlice_l173_253 = (_zz_when_ArraySlice_l173_253_1 <= _zz_when_ArraySlice_l173_253_3);
  assign when_ArraySlice_l165_254 = (_zz_when_ArraySlice_l165_254 <= selectWriteFifo);
  assign when_ArraySlice_l166_254 = (_zz_when_ArraySlice_l166_254 <= _zz_when_ArraySlice_l166_254_2);
  assign _zz_when_ArraySlice_l112_254 = (wReg % _zz__zz_when_ArraySlice_l112_254);
  assign when_ArraySlice_l112_254 = (_zz_when_ArraySlice_l112_254 != 6'h0);
  assign when_ArraySlice_l113_254 = (7'h40 <= _zz_when_ArraySlice_l113_254);
  always @(*) begin
    if(when_ArraySlice_l112_254) begin
      if(when_ArraySlice_l113_254) begin
        _zz_when_ArraySlice_l173_254 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_254 = (_zz__zz_when_ArraySlice_l173_254 - _zz__zz_when_ArraySlice_l173_254_3);
      end
    end else begin
      if(when_ArraySlice_l118_254) begin
        _zz_when_ArraySlice_l173_254 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_254 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_254 = (_zz_when_ArraySlice_l118_254 <= wReg);
  assign when_ArraySlice_l173_254 = (_zz_when_ArraySlice_l173_254_1 <= _zz_when_ArraySlice_l173_254_3);
  assign when_ArraySlice_l165_255 = (_zz_when_ArraySlice_l165_255 <= selectWriteFifo);
  assign when_ArraySlice_l166_255 = (_zz_when_ArraySlice_l166_255 <= _zz_when_ArraySlice_l166_255_2);
  assign _zz_when_ArraySlice_l112_255 = (wReg % _zz__zz_when_ArraySlice_l112_255);
  assign when_ArraySlice_l112_255 = (_zz_when_ArraySlice_l112_255 != 6'h0);
  assign when_ArraySlice_l113_255 = (7'h40 <= _zz_when_ArraySlice_l113_255);
  always @(*) begin
    if(when_ArraySlice_l112_255) begin
      if(when_ArraySlice_l113_255) begin
        _zz_when_ArraySlice_l173_255 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_255 = (_zz__zz_when_ArraySlice_l173_255 - _zz__zz_when_ArraySlice_l173_255_3);
      end
    end else begin
      if(when_ArraySlice_l118_255) begin
        _zz_when_ArraySlice_l173_255 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_255 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_255 = (_zz_when_ArraySlice_l118_255 <= wReg);
  assign when_ArraySlice_l173_255 = (_zz_when_ArraySlice_l173_255_1 <= _zz_when_ArraySlice_l173_255_3);
  assign when_ArraySlice_l311_1 = (! ((((((_zz_when_ArraySlice_l311_1_1 && _zz_when_ArraySlice_l311_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l311_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l311_1_4 && _zz_when_ArraySlice_l311_1_5) && (debug_4_31 == _zz_when_ArraySlice_l311_1_6)) && (debug_5_31 == 1'b1)) && (debug_6_31 == 1'b1)) && (debug_7_31 == 1'b1))));
  assign outputStreamArrayData_1_fire_12 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l315_1 = ((_zz_when_ArraySlice_l315_1_1 == 13'h0) && outputStreamArrayData_1_fire_12);
  assign when_ArraySlice_l301_1 = (allowPadding_1 && (wReg <= _zz_when_ArraySlice_l301_1_1));
  assign outputStreamArrayData_1_fire_13 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l322_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l322_1_1);
  assign when_ArraySlice_l240_2 = (_zz_when_ArraySlice_l240_2_1 < wReg);
  assign when_ArraySlice_l241_2 = ((! holdReadOp_2) && (_zz_when_ArraySlice_l241_2_1 != 7'h0));
  assign _zz_outputStreamArrayData_2_valid_1 = (selectReadFifo_2 + _zz__zz_outputStreamArrayData_2_valid_1_1);
  assign _zz_13 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_2_valid_1);
  assign _zz_io_pop_ready_10 = outputStreamArrayData_2_ready;
  assign when_ArraySlice_l246_2 = (! holdReadOp_2);
  assign outputStreamArrayData_2_fire_7 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l247_2 = ((_zz_when_ArraySlice_l247_2_1 < _zz_when_ArraySlice_l247_2_3) && outputStreamArrayData_2_fire_7);
  assign when_ArraySlice_l248_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l248_2_1);
  assign when_ArraySlice_l251_2 = (_zz_when_ArraySlice_l251_2_1 == 13'h0);
  assign outputStreamArrayData_2_fire_8 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l256_2 = ((_zz_when_ArraySlice_l256_2_1 == _zz_when_ArraySlice_l256_2_5) && outputStreamArrayData_2_fire_8);
  assign when_ArraySlice_l257_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l257_2_1);
  assign _zz_when_ArraySlice_l94_30 = (hReg % _zz__zz_when_ArraySlice_l94_30);
  assign when_ArraySlice_l94_30 = (_zz_when_ArraySlice_l94_30 != 6'h0);
  assign when_ArraySlice_l95_30 = (7'h40 <= _zz_when_ArraySlice_l95_30);
  always @(*) begin
    if(when_ArraySlice_l94_30) begin
      if(when_ArraySlice_l95_30) begin
        _zz_when_ArraySlice_l259_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_2 = (_zz__zz_when_ArraySlice_l259_2_1 - _zz__zz_when_ArraySlice_l259_2_4);
      end
    end else begin
      if(when_ArraySlice_l99_30) begin
        _zz_when_ArraySlice_l259_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_2 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_30 = (_zz_when_ArraySlice_l99_30 <= hReg);
  assign when_ArraySlice_l259_2 = (_zz_when_ArraySlice_l259_2_1 < _zz_when_ArraySlice_l259_2_4);
  always @(*) begin
    debug_0_32 = 1'b0;
    if(when_ArraySlice_l165_256) begin
      if(when_ArraySlice_l166_256) begin
        debug_0_32 = 1'b1;
      end else begin
        debug_0_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_256) begin
        debug_0_32 = 1'b1;
      end else begin
        debug_0_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_32 = 1'b0;
    if(when_ArraySlice_l165_257) begin
      if(when_ArraySlice_l166_257) begin
        debug_1_32 = 1'b1;
      end else begin
        debug_1_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_257) begin
        debug_1_32 = 1'b1;
      end else begin
        debug_1_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_32 = 1'b0;
    if(when_ArraySlice_l165_258) begin
      if(when_ArraySlice_l166_258) begin
        debug_2_32 = 1'b1;
      end else begin
        debug_2_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_258) begin
        debug_2_32 = 1'b1;
      end else begin
        debug_2_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_32 = 1'b0;
    if(when_ArraySlice_l165_259) begin
      if(when_ArraySlice_l166_259) begin
        debug_3_32 = 1'b1;
      end else begin
        debug_3_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_259) begin
        debug_3_32 = 1'b1;
      end else begin
        debug_3_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_32 = 1'b0;
    if(when_ArraySlice_l165_260) begin
      if(when_ArraySlice_l166_260) begin
        debug_4_32 = 1'b1;
      end else begin
        debug_4_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_260) begin
        debug_4_32 = 1'b1;
      end else begin
        debug_4_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_32 = 1'b0;
    if(when_ArraySlice_l165_261) begin
      if(when_ArraySlice_l166_261) begin
        debug_5_32 = 1'b1;
      end else begin
        debug_5_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_261) begin
        debug_5_32 = 1'b1;
      end else begin
        debug_5_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_32 = 1'b0;
    if(when_ArraySlice_l165_262) begin
      if(when_ArraySlice_l166_262) begin
        debug_6_32 = 1'b1;
      end else begin
        debug_6_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_262) begin
        debug_6_32 = 1'b1;
      end else begin
        debug_6_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_32 = 1'b0;
    if(when_ArraySlice_l165_263) begin
      if(when_ArraySlice_l166_263) begin
        debug_7_32 = 1'b1;
      end else begin
        debug_7_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_263) begin
        debug_7_32 = 1'b1;
      end else begin
        debug_7_32 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_256 = (_zz_when_ArraySlice_l165_256 <= selectWriteFifo);
  assign when_ArraySlice_l166_256 = (_zz_when_ArraySlice_l166_256 <= _zz_when_ArraySlice_l166_256_1);
  assign _zz_when_ArraySlice_l112_256 = (wReg % _zz__zz_when_ArraySlice_l112_256);
  assign when_ArraySlice_l112_256 = (_zz_when_ArraySlice_l112_256 != 6'h0);
  assign when_ArraySlice_l113_256 = (7'h40 <= _zz_when_ArraySlice_l113_256);
  always @(*) begin
    if(when_ArraySlice_l112_256) begin
      if(when_ArraySlice_l113_256) begin
        _zz_when_ArraySlice_l173_256 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_256 = (_zz__zz_when_ArraySlice_l173_256 - _zz__zz_when_ArraySlice_l173_256_3);
      end
    end else begin
      if(when_ArraySlice_l118_256) begin
        _zz_when_ArraySlice_l173_256 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_256 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_256 = (_zz_when_ArraySlice_l118_256 <= wReg);
  assign when_ArraySlice_l173_256 = (_zz_when_ArraySlice_l173_256_1 <= _zz_when_ArraySlice_l173_256_2);
  assign when_ArraySlice_l165_257 = (_zz_when_ArraySlice_l165_257 <= selectWriteFifo);
  assign when_ArraySlice_l166_257 = (_zz_when_ArraySlice_l166_257 <= _zz_when_ArraySlice_l166_257_1);
  assign _zz_when_ArraySlice_l112_257 = (wReg % _zz__zz_when_ArraySlice_l112_257);
  assign when_ArraySlice_l112_257 = (_zz_when_ArraySlice_l112_257 != 6'h0);
  assign when_ArraySlice_l113_257 = (7'h40 <= _zz_when_ArraySlice_l113_257);
  always @(*) begin
    if(when_ArraySlice_l112_257) begin
      if(when_ArraySlice_l113_257) begin
        _zz_when_ArraySlice_l173_257 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_257 = (_zz__zz_when_ArraySlice_l173_257 - _zz__zz_when_ArraySlice_l173_257_3);
      end
    end else begin
      if(when_ArraySlice_l118_257) begin
        _zz_when_ArraySlice_l173_257 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_257 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_257 = (_zz_when_ArraySlice_l118_257 <= wReg);
  assign when_ArraySlice_l173_257 = (_zz_when_ArraySlice_l173_257_1 <= _zz_when_ArraySlice_l173_257_3);
  assign when_ArraySlice_l165_258 = (_zz_when_ArraySlice_l165_258 <= selectWriteFifo);
  assign when_ArraySlice_l166_258 = (_zz_when_ArraySlice_l166_258 <= _zz_when_ArraySlice_l166_258_1);
  assign _zz_when_ArraySlice_l112_258 = (wReg % _zz__zz_when_ArraySlice_l112_258);
  assign when_ArraySlice_l112_258 = (_zz_when_ArraySlice_l112_258 != 6'h0);
  assign when_ArraySlice_l113_258 = (7'h40 <= _zz_when_ArraySlice_l113_258);
  always @(*) begin
    if(when_ArraySlice_l112_258) begin
      if(when_ArraySlice_l113_258) begin
        _zz_when_ArraySlice_l173_258 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_258 = (_zz__zz_when_ArraySlice_l173_258 - _zz__zz_when_ArraySlice_l173_258_3);
      end
    end else begin
      if(when_ArraySlice_l118_258) begin
        _zz_when_ArraySlice_l173_258 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_258 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_258 = (_zz_when_ArraySlice_l118_258 <= wReg);
  assign when_ArraySlice_l173_258 = (_zz_when_ArraySlice_l173_258_1 <= _zz_when_ArraySlice_l173_258_3);
  assign when_ArraySlice_l165_259 = (_zz_when_ArraySlice_l165_259 <= selectWriteFifo);
  assign when_ArraySlice_l166_259 = (_zz_when_ArraySlice_l166_259 <= _zz_when_ArraySlice_l166_259_1);
  assign _zz_when_ArraySlice_l112_259 = (wReg % _zz__zz_when_ArraySlice_l112_259);
  assign when_ArraySlice_l112_259 = (_zz_when_ArraySlice_l112_259 != 6'h0);
  assign when_ArraySlice_l113_259 = (7'h40 <= _zz_when_ArraySlice_l113_259);
  always @(*) begin
    if(when_ArraySlice_l112_259) begin
      if(when_ArraySlice_l113_259) begin
        _zz_when_ArraySlice_l173_259 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_259 = (_zz__zz_when_ArraySlice_l173_259 - _zz__zz_when_ArraySlice_l173_259_3);
      end
    end else begin
      if(when_ArraySlice_l118_259) begin
        _zz_when_ArraySlice_l173_259 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_259 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_259 = (_zz_when_ArraySlice_l118_259 <= wReg);
  assign when_ArraySlice_l173_259 = (_zz_when_ArraySlice_l173_259_1 <= _zz_when_ArraySlice_l173_259_3);
  assign when_ArraySlice_l165_260 = (_zz_when_ArraySlice_l165_260 <= selectWriteFifo);
  assign when_ArraySlice_l166_260 = (_zz_when_ArraySlice_l166_260 <= _zz_when_ArraySlice_l166_260_1);
  assign _zz_when_ArraySlice_l112_260 = (wReg % _zz__zz_when_ArraySlice_l112_260);
  assign when_ArraySlice_l112_260 = (_zz_when_ArraySlice_l112_260 != 6'h0);
  assign when_ArraySlice_l113_260 = (7'h40 <= _zz_when_ArraySlice_l113_260);
  always @(*) begin
    if(when_ArraySlice_l112_260) begin
      if(when_ArraySlice_l113_260) begin
        _zz_when_ArraySlice_l173_260 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_260 = (_zz__zz_when_ArraySlice_l173_260 - _zz__zz_when_ArraySlice_l173_260_3);
      end
    end else begin
      if(when_ArraySlice_l118_260) begin
        _zz_when_ArraySlice_l173_260 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_260 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_260 = (_zz_when_ArraySlice_l118_260 <= wReg);
  assign when_ArraySlice_l173_260 = (_zz_when_ArraySlice_l173_260_1 <= _zz_when_ArraySlice_l173_260_3);
  assign when_ArraySlice_l165_261 = (_zz_when_ArraySlice_l165_261 <= selectWriteFifo);
  assign when_ArraySlice_l166_261 = (_zz_when_ArraySlice_l166_261 <= _zz_when_ArraySlice_l166_261_2);
  assign _zz_when_ArraySlice_l112_261 = (wReg % _zz__zz_when_ArraySlice_l112_261);
  assign when_ArraySlice_l112_261 = (_zz_when_ArraySlice_l112_261 != 6'h0);
  assign when_ArraySlice_l113_261 = (7'h40 <= _zz_when_ArraySlice_l113_261);
  always @(*) begin
    if(when_ArraySlice_l112_261) begin
      if(when_ArraySlice_l113_261) begin
        _zz_when_ArraySlice_l173_261 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_261 = (_zz__zz_when_ArraySlice_l173_261 - _zz__zz_when_ArraySlice_l173_261_3);
      end
    end else begin
      if(when_ArraySlice_l118_261) begin
        _zz_when_ArraySlice_l173_261 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_261 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_261 = (_zz_when_ArraySlice_l118_261 <= wReg);
  assign when_ArraySlice_l173_261 = (_zz_when_ArraySlice_l173_261_1 <= _zz_when_ArraySlice_l173_261_3);
  assign when_ArraySlice_l165_262 = (_zz_when_ArraySlice_l165_262 <= selectWriteFifo);
  assign when_ArraySlice_l166_262 = (_zz_when_ArraySlice_l166_262 <= _zz_when_ArraySlice_l166_262_2);
  assign _zz_when_ArraySlice_l112_262 = (wReg % _zz__zz_when_ArraySlice_l112_262);
  assign when_ArraySlice_l112_262 = (_zz_when_ArraySlice_l112_262 != 6'h0);
  assign when_ArraySlice_l113_262 = (7'h40 <= _zz_when_ArraySlice_l113_262);
  always @(*) begin
    if(when_ArraySlice_l112_262) begin
      if(when_ArraySlice_l113_262) begin
        _zz_when_ArraySlice_l173_262 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_262 = (_zz__zz_when_ArraySlice_l173_262 - _zz__zz_when_ArraySlice_l173_262_3);
      end
    end else begin
      if(when_ArraySlice_l118_262) begin
        _zz_when_ArraySlice_l173_262 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_262 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_262 = (_zz_when_ArraySlice_l118_262 <= wReg);
  assign when_ArraySlice_l173_262 = (_zz_when_ArraySlice_l173_262_1 <= _zz_when_ArraySlice_l173_262_3);
  assign when_ArraySlice_l165_263 = (_zz_when_ArraySlice_l165_263 <= selectWriteFifo);
  assign when_ArraySlice_l166_263 = (_zz_when_ArraySlice_l166_263 <= _zz_when_ArraySlice_l166_263_2);
  assign _zz_when_ArraySlice_l112_263 = (wReg % _zz__zz_when_ArraySlice_l112_263);
  assign when_ArraySlice_l112_263 = (_zz_when_ArraySlice_l112_263 != 6'h0);
  assign when_ArraySlice_l113_263 = (7'h40 <= _zz_when_ArraySlice_l113_263);
  always @(*) begin
    if(when_ArraySlice_l112_263) begin
      if(when_ArraySlice_l113_263) begin
        _zz_when_ArraySlice_l173_263 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_263 = (_zz__zz_when_ArraySlice_l173_263 - _zz__zz_when_ArraySlice_l173_263_3);
      end
    end else begin
      if(when_ArraySlice_l118_263) begin
        _zz_when_ArraySlice_l173_263 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_263 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_263 = (_zz_when_ArraySlice_l118_263 <= wReg);
  assign when_ArraySlice_l173_263 = (_zz_when_ArraySlice_l173_263_1 <= _zz_when_ArraySlice_l173_263_3);
  assign when_ArraySlice_l265_2 = (! ((((((_zz_when_ArraySlice_l265_2_1 && _zz_when_ArraySlice_l265_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l265_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l265_2_4 && _zz_when_ArraySlice_l265_2_5) && (debug_4_32 == _zz_when_ArraySlice_l265_2_6)) && (debug_5_32 == 1'b1)) && (debug_6_32 == 1'b1)) && (debug_7_32 == 1'b1))));
  assign when_ArraySlice_l268_2 = (wReg <= _zz_when_ArraySlice_l268_2_1);
  assign when_ArraySlice_l272_2 = (_zz_when_ArraySlice_l272_2_1 == 13'h0);
  assign when_ArraySlice_l276_2 = (_zz_when_ArraySlice_l276_2_1 == 7'h0);
  assign outputStreamArrayData_2_fire_9 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l277_2 = ((handshakeTimes_2_value == _zz_when_ArraySlice_l277_2_1) && outputStreamArrayData_2_fire_9);
  assign _zz_when_ArraySlice_l94_31 = (hReg % _zz__zz_when_ArraySlice_l94_31);
  assign when_ArraySlice_l94_31 = (_zz_when_ArraySlice_l94_31 != 6'h0);
  assign when_ArraySlice_l95_31 = (7'h40 <= _zz_when_ArraySlice_l95_31);
  always @(*) begin
    if(when_ArraySlice_l94_31) begin
      if(when_ArraySlice_l95_31) begin
        _zz_when_ArraySlice_l279_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_2 = (_zz__zz_when_ArraySlice_l279_2_1 - _zz__zz_when_ArraySlice_l279_2_4);
      end
    end else begin
      if(when_ArraySlice_l99_31) begin
        _zz_when_ArraySlice_l279_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_2 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_31 = (_zz_when_ArraySlice_l99_31 <= hReg);
  assign when_ArraySlice_l279_2 = (_zz_when_ArraySlice_l279_2_1 < _zz_when_ArraySlice_l279_2_4);
  always @(*) begin
    debug_0_33 = 1'b0;
    if(when_ArraySlice_l165_264) begin
      if(when_ArraySlice_l166_264) begin
        debug_0_33 = 1'b1;
      end else begin
        debug_0_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_264) begin
        debug_0_33 = 1'b1;
      end else begin
        debug_0_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_33 = 1'b0;
    if(when_ArraySlice_l165_265) begin
      if(when_ArraySlice_l166_265) begin
        debug_1_33 = 1'b1;
      end else begin
        debug_1_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_265) begin
        debug_1_33 = 1'b1;
      end else begin
        debug_1_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_33 = 1'b0;
    if(when_ArraySlice_l165_266) begin
      if(when_ArraySlice_l166_266) begin
        debug_2_33 = 1'b1;
      end else begin
        debug_2_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_266) begin
        debug_2_33 = 1'b1;
      end else begin
        debug_2_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_33 = 1'b0;
    if(when_ArraySlice_l165_267) begin
      if(when_ArraySlice_l166_267) begin
        debug_3_33 = 1'b1;
      end else begin
        debug_3_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_267) begin
        debug_3_33 = 1'b1;
      end else begin
        debug_3_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_33 = 1'b0;
    if(when_ArraySlice_l165_268) begin
      if(when_ArraySlice_l166_268) begin
        debug_4_33 = 1'b1;
      end else begin
        debug_4_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_268) begin
        debug_4_33 = 1'b1;
      end else begin
        debug_4_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_33 = 1'b0;
    if(when_ArraySlice_l165_269) begin
      if(when_ArraySlice_l166_269) begin
        debug_5_33 = 1'b1;
      end else begin
        debug_5_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_269) begin
        debug_5_33 = 1'b1;
      end else begin
        debug_5_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_33 = 1'b0;
    if(when_ArraySlice_l165_270) begin
      if(when_ArraySlice_l166_270) begin
        debug_6_33 = 1'b1;
      end else begin
        debug_6_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_270) begin
        debug_6_33 = 1'b1;
      end else begin
        debug_6_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_33 = 1'b0;
    if(when_ArraySlice_l165_271) begin
      if(when_ArraySlice_l166_271) begin
        debug_7_33 = 1'b1;
      end else begin
        debug_7_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_271) begin
        debug_7_33 = 1'b1;
      end else begin
        debug_7_33 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_264 = (_zz_when_ArraySlice_l165_264 <= selectWriteFifo);
  assign when_ArraySlice_l166_264 = (_zz_when_ArraySlice_l166_264 <= _zz_when_ArraySlice_l166_264_1);
  assign _zz_when_ArraySlice_l112_264 = (wReg % _zz__zz_when_ArraySlice_l112_264);
  assign when_ArraySlice_l112_264 = (_zz_when_ArraySlice_l112_264 != 6'h0);
  assign when_ArraySlice_l113_264 = (7'h40 <= _zz_when_ArraySlice_l113_264);
  always @(*) begin
    if(when_ArraySlice_l112_264) begin
      if(when_ArraySlice_l113_264) begin
        _zz_when_ArraySlice_l173_264 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_264 = (_zz__zz_when_ArraySlice_l173_264 - _zz__zz_when_ArraySlice_l173_264_3);
      end
    end else begin
      if(when_ArraySlice_l118_264) begin
        _zz_when_ArraySlice_l173_264 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_264 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_264 = (_zz_when_ArraySlice_l118_264 <= wReg);
  assign when_ArraySlice_l173_264 = (_zz_when_ArraySlice_l173_264_1 <= _zz_when_ArraySlice_l173_264_2);
  assign when_ArraySlice_l165_265 = (_zz_when_ArraySlice_l165_265 <= selectWriteFifo);
  assign when_ArraySlice_l166_265 = (_zz_when_ArraySlice_l166_265 <= _zz_when_ArraySlice_l166_265_1);
  assign _zz_when_ArraySlice_l112_265 = (wReg % _zz__zz_when_ArraySlice_l112_265);
  assign when_ArraySlice_l112_265 = (_zz_when_ArraySlice_l112_265 != 6'h0);
  assign when_ArraySlice_l113_265 = (7'h40 <= _zz_when_ArraySlice_l113_265);
  always @(*) begin
    if(when_ArraySlice_l112_265) begin
      if(when_ArraySlice_l113_265) begin
        _zz_when_ArraySlice_l173_265 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_265 = (_zz__zz_when_ArraySlice_l173_265 - _zz__zz_when_ArraySlice_l173_265_3);
      end
    end else begin
      if(when_ArraySlice_l118_265) begin
        _zz_when_ArraySlice_l173_265 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_265 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_265 = (_zz_when_ArraySlice_l118_265 <= wReg);
  assign when_ArraySlice_l173_265 = (_zz_when_ArraySlice_l173_265_1 <= _zz_when_ArraySlice_l173_265_3);
  assign when_ArraySlice_l165_266 = (_zz_when_ArraySlice_l165_266 <= selectWriteFifo);
  assign when_ArraySlice_l166_266 = (_zz_when_ArraySlice_l166_266 <= _zz_when_ArraySlice_l166_266_1);
  assign _zz_when_ArraySlice_l112_266 = (wReg % _zz__zz_when_ArraySlice_l112_266);
  assign when_ArraySlice_l112_266 = (_zz_when_ArraySlice_l112_266 != 6'h0);
  assign when_ArraySlice_l113_266 = (7'h40 <= _zz_when_ArraySlice_l113_266);
  always @(*) begin
    if(when_ArraySlice_l112_266) begin
      if(when_ArraySlice_l113_266) begin
        _zz_when_ArraySlice_l173_266 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_266 = (_zz__zz_when_ArraySlice_l173_266 - _zz__zz_when_ArraySlice_l173_266_3);
      end
    end else begin
      if(when_ArraySlice_l118_266) begin
        _zz_when_ArraySlice_l173_266 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_266 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_266 = (_zz_when_ArraySlice_l118_266 <= wReg);
  assign when_ArraySlice_l173_266 = (_zz_when_ArraySlice_l173_266_1 <= _zz_when_ArraySlice_l173_266_3);
  assign when_ArraySlice_l165_267 = (_zz_when_ArraySlice_l165_267 <= selectWriteFifo);
  assign when_ArraySlice_l166_267 = (_zz_when_ArraySlice_l166_267 <= _zz_when_ArraySlice_l166_267_1);
  assign _zz_when_ArraySlice_l112_267 = (wReg % _zz__zz_when_ArraySlice_l112_267);
  assign when_ArraySlice_l112_267 = (_zz_when_ArraySlice_l112_267 != 6'h0);
  assign when_ArraySlice_l113_267 = (7'h40 <= _zz_when_ArraySlice_l113_267);
  always @(*) begin
    if(when_ArraySlice_l112_267) begin
      if(when_ArraySlice_l113_267) begin
        _zz_when_ArraySlice_l173_267 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_267 = (_zz__zz_when_ArraySlice_l173_267 - _zz__zz_when_ArraySlice_l173_267_3);
      end
    end else begin
      if(when_ArraySlice_l118_267) begin
        _zz_when_ArraySlice_l173_267 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_267 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_267 = (_zz_when_ArraySlice_l118_267 <= wReg);
  assign when_ArraySlice_l173_267 = (_zz_when_ArraySlice_l173_267_1 <= _zz_when_ArraySlice_l173_267_3);
  assign when_ArraySlice_l165_268 = (_zz_when_ArraySlice_l165_268 <= selectWriteFifo);
  assign when_ArraySlice_l166_268 = (_zz_when_ArraySlice_l166_268 <= _zz_when_ArraySlice_l166_268_1);
  assign _zz_when_ArraySlice_l112_268 = (wReg % _zz__zz_when_ArraySlice_l112_268);
  assign when_ArraySlice_l112_268 = (_zz_when_ArraySlice_l112_268 != 6'h0);
  assign when_ArraySlice_l113_268 = (7'h40 <= _zz_when_ArraySlice_l113_268);
  always @(*) begin
    if(when_ArraySlice_l112_268) begin
      if(when_ArraySlice_l113_268) begin
        _zz_when_ArraySlice_l173_268 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_268 = (_zz__zz_when_ArraySlice_l173_268 - _zz__zz_when_ArraySlice_l173_268_3);
      end
    end else begin
      if(when_ArraySlice_l118_268) begin
        _zz_when_ArraySlice_l173_268 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_268 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_268 = (_zz_when_ArraySlice_l118_268 <= wReg);
  assign when_ArraySlice_l173_268 = (_zz_when_ArraySlice_l173_268_1 <= _zz_when_ArraySlice_l173_268_3);
  assign when_ArraySlice_l165_269 = (_zz_when_ArraySlice_l165_269 <= selectWriteFifo);
  assign when_ArraySlice_l166_269 = (_zz_when_ArraySlice_l166_269 <= _zz_when_ArraySlice_l166_269_2);
  assign _zz_when_ArraySlice_l112_269 = (wReg % _zz__zz_when_ArraySlice_l112_269);
  assign when_ArraySlice_l112_269 = (_zz_when_ArraySlice_l112_269 != 6'h0);
  assign when_ArraySlice_l113_269 = (7'h40 <= _zz_when_ArraySlice_l113_269);
  always @(*) begin
    if(when_ArraySlice_l112_269) begin
      if(when_ArraySlice_l113_269) begin
        _zz_when_ArraySlice_l173_269 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_269 = (_zz__zz_when_ArraySlice_l173_269 - _zz__zz_when_ArraySlice_l173_269_3);
      end
    end else begin
      if(when_ArraySlice_l118_269) begin
        _zz_when_ArraySlice_l173_269 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_269 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_269 = (_zz_when_ArraySlice_l118_269 <= wReg);
  assign when_ArraySlice_l173_269 = (_zz_when_ArraySlice_l173_269_1 <= _zz_when_ArraySlice_l173_269_3);
  assign when_ArraySlice_l165_270 = (_zz_when_ArraySlice_l165_270 <= selectWriteFifo);
  assign when_ArraySlice_l166_270 = (_zz_when_ArraySlice_l166_270 <= _zz_when_ArraySlice_l166_270_2);
  assign _zz_when_ArraySlice_l112_270 = (wReg % _zz__zz_when_ArraySlice_l112_270);
  assign when_ArraySlice_l112_270 = (_zz_when_ArraySlice_l112_270 != 6'h0);
  assign when_ArraySlice_l113_270 = (7'h40 <= _zz_when_ArraySlice_l113_270);
  always @(*) begin
    if(when_ArraySlice_l112_270) begin
      if(when_ArraySlice_l113_270) begin
        _zz_when_ArraySlice_l173_270 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_270 = (_zz__zz_when_ArraySlice_l173_270 - _zz__zz_when_ArraySlice_l173_270_3);
      end
    end else begin
      if(when_ArraySlice_l118_270) begin
        _zz_when_ArraySlice_l173_270 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_270 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_270 = (_zz_when_ArraySlice_l118_270 <= wReg);
  assign when_ArraySlice_l173_270 = (_zz_when_ArraySlice_l173_270_1 <= _zz_when_ArraySlice_l173_270_3);
  assign when_ArraySlice_l165_271 = (_zz_when_ArraySlice_l165_271 <= selectWriteFifo);
  assign when_ArraySlice_l166_271 = (_zz_when_ArraySlice_l166_271 <= _zz_when_ArraySlice_l166_271_2);
  assign _zz_when_ArraySlice_l112_271 = (wReg % _zz__zz_when_ArraySlice_l112_271);
  assign when_ArraySlice_l112_271 = (_zz_when_ArraySlice_l112_271 != 6'h0);
  assign when_ArraySlice_l113_271 = (7'h40 <= _zz_when_ArraySlice_l113_271);
  always @(*) begin
    if(when_ArraySlice_l112_271) begin
      if(when_ArraySlice_l113_271) begin
        _zz_when_ArraySlice_l173_271 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_271 = (_zz__zz_when_ArraySlice_l173_271 - _zz__zz_when_ArraySlice_l173_271_3);
      end
    end else begin
      if(when_ArraySlice_l118_271) begin
        _zz_when_ArraySlice_l173_271 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_271 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_271 = (_zz_when_ArraySlice_l118_271 <= wReg);
  assign when_ArraySlice_l173_271 = (_zz_when_ArraySlice_l173_271_1 <= _zz_when_ArraySlice_l173_271_3);
  assign when_ArraySlice_l285_2 = (! ((((((_zz_when_ArraySlice_l285_2_1 && _zz_when_ArraySlice_l285_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l285_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l285_2_4 && _zz_when_ArraySlice_l285_2_5) && (debug_4_33 == _zz_when_ArraySlice_l285_2_6)) && (debug_5_33 == 1'b1)) && (debug_6_33 == 1'b1)) && (debug_7_33 == 1'b1))));
  assign when_ArraySlice_l288_2 = (wReg <= _zz_when_ArraySlice_l288_2_1);
  assign outputStreamArrayData_2_fire_10 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l292_2 = ((_zz_when_ArraySlice_l292_2_1 == 13'h0) && outputStreamArrayData_2_fire_10);
  assign outputStreamArrayData_2_fire_11 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l303_2 = ((handshakeTimes_2_value == _zz_when_ArraySlice_l303_2_1) && outputStreamArrayData_2_fire_11);
  assign _zz_when_ArraySlice_l94_32 = (hReg % _zz__zz_when_ArraySlice_l94_32);
  assign when_ArraySlice_l94_32 = (_zz_when_ArraySlice_l94_32 != 6'h0);
  assign when_ArraySlice_l95_32 = (7'h40 <= _zz_when_ArraySlice_l95_32);
  always @(*) begin
    if(when_ArraySlice_l94_32) begin
      if(when_ArraySlice_l95_32) begin
        _zz_when_ArraySlice_l304_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_2 = (_zz__zz_when_ArraySlice_l304_2_1 - _zz__zz_when_ArraySlice_l304_2_4);
      end
    end else begin
      if(when_ArraySlice_l99_32) begin
        _zz_when_ArraySlice_l304_2 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_2 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_32 = (_zz_when_ArraySlice_l99_32 <= hReg);
  assign when_ArraySlice_l304_2 = (_zz_when_ArraySlice_l304_2_1 < _zz_when_ArraySlice_l304_2_4);
  always @(*) begin
    debug_0_34 = 1'b0;
    if(when_ArraySlice_l165_272) begin
      if(when_ArraySlice_l166_272) begin
        debug_0_34 = 1'b1;
      end else begin
        debug_0_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_272) begin
        debug_0_34 = 1'b1;
      end else begin
        debug_0_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_34 = 1'b0;
    if(when_ArraySlice_l165_273) begin
      if(when_ArraySlice_l166_273) begin
        debug_1_34 = 1'b1;
      end else begin
        debug_1_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_273) begin
        debug_1_34 = 1'b1;
      end else begin
        debug_1_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_34 = 1'b0;
    if(when_ArraySlice_l165_274) begin
      if(when_ArraySlice_l166_274) begin
        debug_2_34 = 1'b1;
      end else begin
        debug_2_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_274) begin
        debug_2_34 = 1'b1;
      end else begin
        debug_2_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_34 = 1'b0;
    if(when_ArraySlice_l165_275) begin
      if(when_ArraySlice_l166_275) begin
        debug_3_34 = 1'b1;
      end else begin
        debug_3_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_275) begin
        debug_3_34 = 1'b1;
      end else begin
        debug_3_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_34 = 1'b0;
    if(when_ArraySlice_l165_276) begin
      if(when_ArraySlice_l166_276) begin
        debug_4_34 = 1'b1;
      end else begin
        debug_4_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_276) begin
        debug_4_34 = 1'b1;
      end else begin
        debug_4_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_34 = 1'b0;
    if(when_ArraySlice_l165_277) begin
      if(when_ArraySlice_l166_277) begin
        debug_5_34 = 1'b1;
      end else begin
        debug_5_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_277) begin
        debug_5_34 = 1'b1;
      end else begin
        debug_5_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_34 = 1'b0;
    if(when_ArraySlice_l165_278) begin
      if(when_ArraySlice_l166_278) begin
        debug_6_34 = 1'b1;
      end else begin
        debug_6_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_278) begin
        debug_6_34 = 1'b1;
      end else begin
        debug_6_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_34 = 1'b0;
    if(when_ArraySlice_l165_279) begin
      if(when_ArraySlice_l166_279) begin
        debug_7_34 = 1'b1;
      end else begin
        debug_7_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_279) begin
        debug_7_34 = 1'b1;
      end else begin
        debug_7_34 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_272 = (_zz_when_ArraySlice_l165_272 <= selectWriteFifo);
  assign when_ArraySlice_l166_272 = (_zz_when_ArraySlice_l166_272 <= _zz_when_ArraySlice_l166_272_1);
  assign _zz_when_ArraySlice_l112_272 = (wReg % _zz__zz_when_ArraySlice_l112_272);
  assign when_ArraySlice_l112_272 = (_zz_when_ArraySlice_l112_272 != 6'h0);
  assign when_ArraySlice_l113_272 = (7'h40 <= _zz_when_ArraySlice_l113_272);
  always @(*) begin
    if(when_ArraySlice_l112_272) begin
      if(when_ArraySlice_l113_272) begin
        _zz_when_ArraySlice_l173_272 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_272 = (_zz__zz_when_ArraySlice_l173_272 - _zz__zz_when_ArraySlice_l173_272_3);
      end
    end else begin
      if(when_ArraySlice_l118_272) begin
        _zz_when_ArraySlice_l173_272 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_272 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_272 = (_zz_when_ArraySlice_l118_272 <= wReg);
  assign when_ArraySlice_l173_272 = (_zz_when_ArraySlice_l173_272_1 <= _zz_when_ArraySlice_l173_272_2);
  assign when_ArraySlice_l165_273 = (_zz_when_ArraySlice_l165_273 <= selectWriteFifo);
  assign when_ArraySlice_l166_273 = (_zz_when_ArraySlice_l166_273 <= _zz_when_ArraySlice_l166_273_1);
  assign _zz_when_ArraySlice_l112_273 = (wReg % _zz__zz_when_ArraySlice_l112_273);
  assign when_ArraySlice_l112_273 = (_zz_when_ArraySlice_l112_273 != 6'h0);
  assign when_ArraySlice_l113_273 = (7'h40 <= _zz_when_ArraySlice_l113_273);
  always @(*) begin
    if(when_ArraySlice_l112_273) begin
      if(when_ArraySlice_l113_273) begin
        _zz_when_ArraySlice_l173_273 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_273 = (_zz__zz_when_ArraySlice_l173_273 - _zz__zz_when_ArraySlice_l173_273_3);
      end
    end else begin
      if(when_ArraySlice_l118_273) begin
        _zz_when_ArraySlice_l173_273 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_273 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_273 = (_zz_when_ArraySlice_l118_273 <= wReg);
  assign when_ArraySlice_l173_273 = (_zz_when_ArraySlice_l173_273_1 <= _zz_when_ArraySlice_l173_273_3);
  assign when_ArraySlice_l165_274 = (_zz_when_ArraySlice_l165_274 <= selectWriteFifo);
  assign when_ArraySlice_l166_274 = (_zz_when_ArraySlice_l166_274 <= _zz_when_ArraySlice_l166_274_1);
  assign _zz_when_ArraySlice_l112_274 = (wReg % _zz__zz_when_ArraySlice_l112_274);
  assign when_ArraySlice_l112_274 = (_zz_when_ArraySlice_l112_274 != 6'h0);
  assign when_ArraySlice_l113_274 = (7'h40 <= _zz_when_ArraySlice_l113_274);
  always @(*) begin
    if(when_ArraySlice_l112_274) begin
      if(when_ArraySlice_l113_274) begin
        _zz_when_ArraySlice_l173_274 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_274 = (_zz__zz_when_ArraySlice_l173_274 - _zz__zz_when_ArraySlice_l173_274_3);
      end
    end else begin
      if(when_ArraySlice_l118_274) begin
        _zz_when_ArraySlice_l173_274 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_274 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_274 = (_zz_when_ArraySlice_l118_274 <= wReg);
  assign when_ArraySlice_l173_274 = (_zz_when_ArraySlice_l173_274_1 <= _zz_when_ArraySlice_l173_274_3);
  assign when_ArraySlice_l165_275 = (_zz_when_ArraySlice_l165_275 <= selectWriteFifo);
  assign when_ArraySlice_l166_275 = (_zz_when_ArraySlice_l166_275 <= _zz_when_ArraySlice_l166_275_1);
  assign _zz_when_ArraySlice_l112_275 = (wReg % _zz__zz_when_ArraySlice_l112_275);
  assign when_ArraySlice_l112_275 = (_zz_when_ArraySlice_l112_275 != 6'h0);
  assign when_ArraySlice_l113_275 = (7'h40 <= _zz_when_ArraySlice_l113_275);
  always @(*) begin
    if(when_ArraySlice_l112_275) begin
      if(when_ArraySlice_l113_275) begin
        _zz_when_ArraySlice_l173_275 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_275 = (_zz__zz_when_ArraySlice_l173_275 - _zz__zz_when_ArraySlice_l173_275_3);
      end
    end else begin
      if(when_ArraySlice_l118_275) begin
        _zz_when_ArraySlice_l173_275 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_275 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_275 = (_zz_when_ArraySlice_l118_275 <= wReg);
  assign when_ArraySlice_l173_275 = (_zz_when_ArraySlice_l173_275_1 <= _zz_when_ArraySlice_l173_275_3);
  assign when_ArraySlice_l165_276 = (_zz_when_ArraySlice_l165_276 <= selectWriteFifo);
  assign when_ArraySlice_l166_276 = (_zz_when_ArraySlice_l166_276 <= _zz_when_ArraySlice_l166_276_1);
  assign _zz_when_ArraySlice_l112_276 = (wReg % _zz__zz_when_ArraySlice_l112_276);
  assign when_ArraySlice_l112_276 = (_zz_when_ArraySlice_l112_276 != 6'h0);
  assign when_ArraySlice_l113_276 = (7'h40 <= _zz_when_ArraySlice_l113_276);
  always @(*) begin
    if(when_ArraySlice_l112_276) begin
      if(when_ArraySlice_l113_276) begin
        _zz_when_ArraySlice_l173_276 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_276 = (_zz__zz_when_ArraySlice_l173_276 - _zz__zz_when_ArraySlice_l173_276_3);
      end
    end else begin
      if(when_ArraySlice_l118_276) begin
        _zz_when_ArraySlice_l173_276 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_276 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_276 = (_zz_when_ArraySlice_l118_276 <= wReg);
  assign when_ArraySlice_l173_276 = (_zz_when_ArraySlice_l173_276_1 <= _zz_when_ArraySlice_l173_276_3);
  assign when_ArraySlice_l165_277 = (_zz_when_ArraySlice_l165_277 <= selectWriteFifo);
  assign when_ArraySlice_l166_277 = (_zz_when_ArraySlice_l166_277 <= _zz_when_ArraySlice_l166_277_2);
  assign _zz_when_ArraySlice_l112_277 = (wReg % _zz__zz_when_ArraySlice_l112_277);
  assign when_ArraySlice_l112_277 = (_zz_when_ArraySlice_l112_277 != 6'h0);
  assign when_ArraySlice_l113_277 = (7'h40 <= _zz_when_ArraySlice_l113_277);
  always @(*) begin
    if(when_ArraySlice_l112_277) begin
      if(when_ArraySlice_l113_277) begin
        _zz_when_ArraySlice_l173_277 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_277 = (_zz__zz_when_ArraySlice_l173_277 - _zz__zz_when_ArraySlice_l173_277_3);
      end
    end else begin
      if(when_ArraySlice_l118_277) begin
        _zz_when_ArraySlice_l173_277 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_277 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_277 = (_zz_when_ArraySlice_l118_277 <= wReg);
  assign when_ArraySlice_l173_277 = (_zz_when_ArraySlice_l173_277_1 <= _zz_when_ArraySlice_l173_277_3);
  assign when_ArraySlice_l165_278 = (_zz_when_ArraySlice_l165_278 <= selectWriteFifo);
  assign when_ArraySlice_l166_278 = (_zz_when_ArraySlice_l166_278 <= _zz_when_ArraySlice_l166_278_2);
  assign _zz_when_ArraySlice_l112_278 = (wReg % _zz__zz_when_ArraySlice_l112_278);
  assign when_ArraySlice_l112_278 = (_zz_when_ArraySlice_l112_278 != 6'h0);
  assign when_ArraySlice_l113_278 = (7'h40 <= _zz_when_ArraySlice_l113_278);
  always @(*) begin
    if(when_ArraySlice_l112_278) begin
      if(when_ArraySlice_l113_278) begin
        _zz_when_ArraySlice_l173_278 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_278 = (_zz__zz_when_ArraySlice_l173_278 - _zz__zz_when_ArraySlice_l173_278_3);
      end
    end else begin
      if(when_ArraySlice_l118_278) begin
        _zz_when_ArraySlice_l173_278 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_278 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_278 = (_zz_when_ArraySlice_l118_278 <= wReg);
  assign when_ArraySlice_l173_278 = (_zz_when_ArraySlice_l173_278_1 <= _zz_when_ArraySlice_l173_278_3);
  assign when_ArraySlice_l165_279 = (_zz_when_ArraySlice_l165_279 <= selectWriteFifo);
  assign when_ArraySlice_l166_279 = (_zz_when_ArraySlice_l166_279 <= _zz_when_ArraySlice_l166_279_2);
  assign _zz_when_ArraySlice_l112_279 = (wReg % _zz__zz_when_ArraySlice_l112_279);
  assign when_ArraySlice_l112_279 = (_zz_when_ArraySlice_l112_279 != 6'h0);
  assign when_ArraySlice_l113_279 = (7'h40 <= _zz_when_ArraySlice_l113_279);
  always @(*) begin
    if(when_ArraySlice_l112_279) begin
      if(when_ArraySlice_l113_279) begin
        _zz_when_ArraySlice_l173_279 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_279 = (_zz__zz_when_ArraySlice_l173_279 - _zz__zz_when_ArraySlice_l173_279_3);
      end
    end else begin
      if(when_ArraySlice_l118_279) begin
        _zz_when_ArraySlice_l173_279 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_279 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_279 = (_zz_when_ArraySlice_l118_279 <= wReg);
  assign when_ArraySlice_l173_279 = (_zz_when_ArraySlice_l173_279_1 <= _zz_when_ArraySlice_l173_279_3);
  assign when_ArraySlice_l311_2 = (! ((((((_zz_when_ArraySlice_l311_2_1 && _zz_when_ArraySlice_l311_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l311_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l311_2_4 && _zz_when_ArraySlice_l311_2_5) && (debug_4_34 == _zz_when_ArraySlice_l311_2_6)) && (debug_5_34 == 1'b1)) && (debug_6_34 == 1'b1)) && (debug_7_34 == 1'b1))));
  assign outputStreamArrayData_2_fire_12 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l315_2 = ((_zz_when_ArraySlice_l315_2_1 == 13'h0) && outputStreamArrayData_2_fire_12);
  assign when_ArraySlice_l301_2 = (allowPadding_2 && (wReg <= _zz_when_ArraySlice_l301_2_1));
  assign outputStreamArrayData_2_fire_13 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l322_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l322_2_1);
  assign when_ArraySlice_l240_3 = (_zz_when_ArraySlice_l240_3 < wReg);
  assign when_ArraySlice_l241_3 = ((! holdReadOp_3) && (_zz_when_ArraySlice_l241_3_1 != 7'h0));
  assign _zz_outputStreamArrayData_3_valid_1 = (selectReadFifo_3 + _zz__zz_outputStreamArrayData_3_valid_1_1);
  assign _zz_14 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_3_valid_1);
  assign _zz_io_pop_ready_11 = outputStreamArrayData_3_ready;
  assign when_ArraySlice_l246_3 = (! holdReadOp_3);
  assign outputStreamArrayData_3_fire_7 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l247_3 = ((_zz_when_ArraySlice_l247_3_1 < _zz_when_ArraySlice_l247_3_3) && outputStreamArrayData_3_fire_7);
  assign when_ArraySlice_l248_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l248_3_1);
  assign when_ArraySlice_l251_3 = (_zz_when_ArraySlice_l251_3_1 == 13'h0);
  assign outputStreamArrayData_3_fire_8 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l256_3 = ((_zz_when_ArraySlice_l256_3_1 == _zz_when_ArraySlice_l256_3_5) && outputStreamArrayData_3_fire_8);
  assign when_ArraySlice_l257_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l257_3_1);
  assign _zz_when_ArraySlice_l94_33 = (hReg % _zz__zz_when_ArraySlice_l94_33);
  assign when_ArraySlice_l94_33 = (_zz_when_ArraySlice_l94_33 != 6'h0);
  assign when_ArraySlice_l95_33 = (7'h40 <= _zz_when_ArraySlice_l95_33);
  always @(*) begin
    if(when_ArraySlice_l94_33) begin
      if(when_ArraySlice_l95_33) begin
        _zz_when_ArraySlice_l259_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_3 = (_zz__zz_when_ArraySlice_l259_3_1 - _zz__zz_when_ArraySlice_l259_3_4);
      end
    end else begin
      if(when_ArraySlice_l99_33) begin
        _zz_when_ArraySlice_l259_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_3 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_33 = (_zz_when_ArraySlice_l99_33 <= hReg);
  assign when_ArraySlice_l259_3 = (_zz_when_ArraySlice_l259_3_1 < _zz_when_ArraySlice_l259_3_4);
  always @(*) begin
    debug_0_35 = 1'b0;
    if(when_ArraySlice_l165_280) begin
      if(when_ArraySlice_l166_280) begin
        debug_0_35 = 1'b1;
      end else begin
        debug_0_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_280) begin
        debug_0_35 = 1'b1;
      end else begin
        debug_0_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_35 = 1'b0;
    if(when_ArraySlice_l165_281) begin
      if(when_ArraySlice_l166_281) begin
        debug_1_35 = 1'b1;
      end else begin
        debug_1_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_281) begin
        debug_1_35 = 1'b1;
      end else begin
        debug_1_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_35 = 1'b0;
    if(when_ArraySlice_l165_282) begin
      if(when_ArraySlice_l166_282) begin
        debug_2_35 = 1'b1;
      end else begin
        debug_2_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_282) begin
        debug_2_35 = 1'b1;
      end else begin
        debug_2_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_35 = 1'b0;
    if(when_ArraySlice_l165_283) begin
      if(when_ArraySlice_l166_283) begin
        debug_3_35 = 1'b1;
      end else begin
        debug_3_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_283) begin
        debug_3_35 = 1'b1;
      end else begin
        debug_3_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_35 = 1'b0;
    if(when_ArraySlice_l165_284) begin
      if(when_ArraySlice_l166_284) begin
        debug_4_35 = 1'b1;
      end else begin
        debug_4_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_284) begin
        debug_4_35 = 1'b1;
      end else begin
        debug_4_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_35 = 1'b0;
    if(when_ArraySlice_l165_285) begin
      if(when_ArraySlice_l166_285) begin
        debug_5_35 = 1'b1;
      end else begin
        debug_5_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_285) begin
        debug_5_35 = 1'b1;
      end else begin
        debug_5_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_35 = 1'b0;
    if(when_ArraySlice_l165_286) begin
      if(when_ArraySlice_l166_286) begin
        debug_6_35 = 1'b1;
      end else begin
        debug_6_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_286) begin
        debug_6_35 = 1'b1;
      end else begin
        debug_6_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_35 = 1'b0;
    if(when_ArraySlice_l165_287) begin
      if(when_ArraySlice_l166_287) begin
        debug_7_35 = 1'b1;
      end else begin
        debug_7_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_287) begin
        debug_7_35 = 1'b1;
      end else begin
        debug_7_35 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_280 = (_zz_when_ArraySlice_l165_280 <= selectWriteFifo);
  assign when_ArraySlice_l166_280 = (_zz_when_ArraySlice_l166_280 <= _zz_when_ArraySlice_l166_280_1);
  assign _zz_when_ArraySlice_l112_280 = (wReg % _zz__zz_when_ArraySlice_l112_280);
  assign when_ArraySlice_l112_280 = (_zz_when_ArraySlice_l112_280 != 6'h0);
  assign when_ArraySlice_l113_280 = (7'h40 <= _zz_when_ArraySlice_l113_280);
  always @(*) begin
    if(when_ArraySlice_l112_280) begin
      if(when_ArraySlice_l113_280) begin
        _zz_when_ArraySlice_l173_280 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_280 = (_zz__zz_when_ArraySlice_l173_280 - _zz__zz_when_ArraySlice_l173_280_3);
      end
    end else begin
      if(when_ArraySlice_l118_280) begin
        _zz_when_ArraySlice_l173_280 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_280 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_280 = (_zz_when_ArraySlice_l118_280 <= wReg);
  assign when_ArraySlice_l173_280 = (_zz_when_ArraySlice_l173_280_1 <= _zz_when_ArraySlice_l173_280_2);
  assign when_ArraySlice_l165_281 = (_zz_when_ArraySlice_l165_281 <= selectWriteFifo);
  assign when_ArraySlice_l166_281 = (_zz_when_ArraySlice_l166_281 <= _zz_when_ArraySlice_l166_281_1);
  assign _zz_when_ArraySlice_l112_281 = (wReg % _zz__zz_when_ArraySlice_l112_281);
  assign when_ArraySlice_l112_281 = (_zz_when_ArraySlice_l112_281 != 6'h0);
  assign when_ArraySlice_l113_281 = (7'h40 <= _zz_when_ArraySlice_l113_281);
  always @(*) begin
    if(when_ArraySlice_l112_281) begin
      if(when_ArraySlice_l113_281) begin
        _zz_when_ArraySlice_l173_281 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_281 = (_zz__zz_when_ArraySlice_l173_281 - _zz__zz_when_ArraySlice_l173_281_3);
      end
    end else begin
      if(when_ArraySlice_l118_281) begin
        _zz_when_ArraySlice_l173_281 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_281 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_281 = (_zz_when_ArraySlice_l118_281 <= wReg);
  assign when_ArraySlice_l173_281 = (_zz_when_ArraySlice_l173_281_1 <= _zz_when_ArraySlice_l173_281_3);
  assign when_ArraySlice_l165_282 = (_zz_when_ArraySlice_l165_282 <= selectWriteFifo);
  assign when_ArraySlice_l166_282 = (_zz_when_ArraySlice_l166_282 <= _zz_when_ArraySlice_l166_282_1);
  assign _zz_when_ArraySlice_l112_282 = (wReg % _zz__zz_when_ArraySlice_l112_282);
  assign when_ArraySlice_l112_282 = (_zz_when_ArraySlice_l112_282 != 6'h0);
  assign when_ArraySlice_l113_282 = (7'h40 <= _zz_when_ArraySlice_l113_282);
  always @(*) begin
    if(when_ArraySlice_l112_282) begin
      if(when_ArraySlice_l113_282) begin
        _zz_when_ArraySlice_l173_282 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_282 = (_zz__zz_when_ArraySlice_l173_282 - _zz__zz_when_ArraySlice_l173_282_3);
      end
    end else begin
      if(when_ArraySlice_l118_282) begin
        _zz_when_ArraySlice_l173_282 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_282 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_282 = (_zz_when_ArraySlice_l118_282 <= wReg);
  assign when_ArraySlice_l173_282 = (_zz_when_ArraySlice_l173_282_1 <= _zz_when_ArraySlice_l173_282_3);
  assign when_ArraySlice_l165_283 = (_zz_when_ArraySlice_l165_283 <= selectWriteFifo);
  assign when_ArraySlice_l166_283 = (_zz_when_ArraySlice_l166_283 <= _zz_when_ArraySlice_l166_283_1);
  assign _zz_when_ArraySlice_l112_283 = (wReg % _zz__zz_when_ArraySlice_l112_283);
  assign when_ArraySlice_l112_283 = (_zz_when_ArraySlice_l112_283 != 6'h0);
  assign when_ArraySlice_l113_283 = (7'h40 <= _zz_when_ArraySlice_l113_283);
  always @(*) begin
    if(when_ArraySlice_l112_283) begin
      if(when_ArraySlice_l113_283) begin
        _zz_when_ArraySlice_l173_283 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_283 = (_zz__zz_when_ArraySlice_l173_283 - _zz__zz_when_ArraySlice_l173_283_3);
      end
    end else begin
      if(when_ArraySlice_l118_283) begin
        _zz_when_ArraySlice_l173_283 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_283 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_283 = (_zz_when_ArraySlice_l118_283 <= wReg);
  assign when_ArraySlice_l173_283 = (_zz_when_ArraySlice_l173_283_1 <= _zz_when_ArraySlice_l173_283_3);
  assign when_ArraySlice_l165_284 = (_zz_when_ArraySlice_l165_284 <= selectWriteFifo);
  assign when_ArraySlice_l166_284 = (_zz_when_ArraySlice_l166_284 <= _zz_when_ArraySlice_l166_284_1);
  assign _zz_when_ArraySlice_l112_284 = (wReg % _zz__zz_when_ArraySlice_l112_284);
  assign when_ArraySlice_l112_284 = (_zz_when_ArraySlice_l112_284 != 6'h0);
  assign when_ArraySlice_l113_284 = (7'h40 <= _zz_when_ArraySlice_l113_284);
  always @(*) begin
    if(when_ArraySlice_l112_284) begin
      if(when_ArraySlice_l113_284) begin
        _zz_when_ArraySlice_l173_284 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_284 = (_zz__zz_when_ArraySlice_l173_284 - _zz__zz_when_ArraySlice_l173_284_3);
      end
    end else begin
      if(when_ArraySlice_l118_284) begin
        _zz_when_ArraySlice_l173_284 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_284 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_284 = (_zz_when_ArraySlice_l118_284 <= wReg);
  assign when_ArraySlice_l173_284 = (_zz_when_ArraySlice_l173_284_1 <= _zz_when_ArraySlice_l173_284_3);
  assign when_ArraySlice_l165_285 = (_zz_when_ArraySlice_l165_285 <= selectWriteFifo);
  assign when_ArraySlice_l166_285 = (_zz_when_ArraySlice_l166_285 <= _zz_when_ArraySlice_l166_285_2);
  assign _zz_when_ArraySlice_l112_285 = (wReg % _zz__zz_when_ArraySlice_l112_285);
  assign when_ArraySlice_l112_285 = (_zz_when_ArraySlice_l112_285 != 6'h0);
  assign when_ArraySlice_l113_285 = (7'h40 <= _zz_when_ArraySlice_l113_285);
  always @(*) begin
    if(when_ArraySlice_l112_285) begin
      if(when_ArraySlice_l113_285) begin
        _zz_when_ArraySlice_l173_285 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_285 = (_zz__zz_when_ArraySlice_l173_285 - _zz__zz_when_ArraySlice_l173_285_3);
      end
    end else begin
      if(when_ArraySlice_l118_285) begin
        _zz_when_ArraySlice_l173_285 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_285 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_285 = (_zz_when_ArraySlice_l118_285 <= wReg);
  assign when_ArraySlice_l173_285 = (_zz_when_ArraySlice_l173_285_1 <= _zz_when_ArraySlice_l173_285_3);
  assign when_ArraySlice_l165_286 = (_zz_when_ArraySlice_l165_286 <= selectWriteFifo);
  assign when_ArraySlice_l166_286 = (_zz_when_ArraySlice_l166_286 <= _zz_when_ArraySlice_l166_286_2);
  assign _zz_when_ArraySlice_l112_286 = (wReg % _zz__zz_when_ArraySlice_l112_286);
  assign when_ArraySlice_l112_286 = (_zz_when_ArraySlice_l112_286 != 6'h0);
  assign when_ArraySlice_l113_286 = (7'h40 <= _zz_when_ArraySlice_l113_286);
  always @(*) begin
    if(when_ArraySlice_l112_286) begin
      if(when_ArraySlice_l113_286) begin
        _zz_when_ArraySlice_l173_286 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_286 = (_zz__zz_when_ArraySlice_l173_286 - _zz__zz_when_ArraySlice_l173_286_3);
      end
    end else begin
      if(when_ArraySlice_l118_286) begin
        _zz_when_ArraySlice_l173_286 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_286 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_286 = (_zz_when_ArraySlice_l118_286 <= wReg);
  assign when_ArraySlice_l173_286 = (_zz_when_ArraySlice_l173_286_1 <= _zz_when_ArraySlice_l173_286_3);
  assign when_ArraySlice_l165_287 = (_zz_when_ArraySlice_l165_287 <= selectWriteFifo);
  assign when_ArraySlice_l166_287 = (_zz_when_ArraySlice_l166_287 <= _zz_when_ArraySlice_l166_287_2);
  assign _zz_when_ArraySlice_l112_287 = (wReg % _zz__zz_when_ArraySlice_l112_287);
  assign when_ArraySlice_l112_287 = (_zz_when_ArraySlice_l112_287 != 6'h0);
  assign when_ArraySlice_l113_287 = (7'h40 <= _zz_when_ArraySlice_l113_287);
  always @(*) begin
    if(when_ArraySlice_l112_287) begin
      if(when_ArraySlice_l113_287) begin
        _zz_when_ArraySlice_l173_287 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_287 = (_zz__zz_when_ArraySlice_l173_287 - _zz__zz_when_ArraySlice_l173_287_3);
      end
    end else begin
      if(when_ArraySlice_l118_287) begin
        _zz_when_ArraySlice_l173_287 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_287 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_287 = (_zz_when_ArraySlice_l118_287 <= wReg);
  assign when_ArraySlice_l173_287 = (_zz_when_ArraySlice_l173_287_1 <= _zz_when_ArraySlice_l173_287_3);
  assign when_ArraySlice_l265_3 = (! ((((((_zz_when_ArraySlice_l265_3_1 && _zz_when_ArraySlice_l265_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l265_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l265_3_4 && _zz_when_ArraySlice_l265_3_5) && (debug_4_35 == _zz_when_ArraySlice_l265_3_6)) && (debug_5_35 == 1'b1)) && (debug_6_35 == 1'b1)) && (debug_7_35 == 1'b1))));
  assign when_ArraySlice_l268_3 = (wReg <= _zz_when_ArraySlice_l268_3_1);
  assign when_ArraySlice_l272_3 = (_zz_when_ArraySlice_l272_3_1 == 13'h0);
  assign when_ArraySlice_l276_3 = (_zz_when_ArraySlice_l276_3_1 == 7'h0);
  assign outputStreamArrayData_3_fire_9 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l277_3 = ((handshakeTimes_3_value == _zz_when_ArraySlice_l277_3_1) && outputStreamArrayData_3_fire_9);
  assign _zz_when_ArraySlice_l94_34 = (hReg % _zz__zz_when_ArraySlice_l94_34);
  assign when_ArraySlice_l94_34 = (_zz_when_ArraySlice_l94_34 != 6'h0);
  assign when_ArraySlice_l95_34 = (7'h40 <= _zz_when_ArraySlice_l95_34);
  always @(*) begin
    if(when_ArraySlice_l94_34) begin
      if(when_ArraySlice_l95_34) begin
        _zz_when_ArraySlice_l279_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_3 = (_zz__zz_when_ArraySlice_l279_3_1 - _zz__zz_when_ArraySlice_l279_3_4);
      end
    end else begin
      if(when_ArraySlice_l99_34) begin
        _zz_when_ArraySlice_l279_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_3 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_34 = (_zz_when_ArraySlice_l99_34 <= hReg);
  assign when_ArraySlice_l279_3 = (_zz_when_ArraySlice_l279_3_1 < _zz_when_ArraySlice_l279_3_4);
  always @(*) begin
    debug_0_36 = 1'b0;
    if(when_ArraySlice_l165_288) begin
      if(when_ArraySlice_l166_288) begin
        debug_0_36 = 1'b1;
      end else begin
        debug_0_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_288) begin
        debug_0_36 = 1'b1;
      end else begin
        debug_0_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_36 = 1'b0;
    if(when_ArraySlice_l165_289) begin
      if(when_ArraySlice_l166_289) begin
        debug_1_36 = 1'b1;
      end else begin
        debug_1_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_289) begin
        debug_1_36 = 1'b1;
      end else begin
        debug_1_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_36 = 1'b0;
    if(when_ArraySlice_l165_290) begin
      if(when_ArraySlice_l166_290) begin
        debug_2_36 = 1'b1;
      end else begin
        debug_2_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_290) begin
        debug_2_36 = 1'b1;
      end else begin
        debug_2_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_36 = 1'b0;
    if(when_ArraySlice_l165_291) begin
      if(when_ArraySlice_l166_291) begin
        debug_3_36 = 1'b1;
      end else begin
        debug_3_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_291) begin
        debug_3_36 = 1'b1;
      end else begin
        debug_3_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_36 = 1'b0;
    if(when_ArraySlice_l165_292) begin
      if(when_ArraySlice_l166_292) begin
        debug_4_36 = 1'b1;
      end else begin
        debug_4_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_292) begin
        debug_4_36 = 1'b1;
      end else begin
        debug_4_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_36 = 1'b0;
    if(when_ArraySlice_l165_293) begin
      if(when_ArraySlice_l166_293) begin
        debug_5_36 = 1'b1;
      end else begin
        debug_5_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_293) begin
        debug_5_36 = 1'b1;
      end else begin
        debug_5_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_36 = 1'b0;
    if(when_ArraySlice_l165_294) begin
      if(when_ArraySlice_l166_294) begin
        debug_6_36 = 1'b1;
      end else begin
        debug_6_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_294) begin
        debug_6_36 = 1'b1;
      end else begin
        debug_6_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_36 = 1'b0;
    if(when_ArraySlice_l165_295) begin
      if(when_ArraySlice_l166_295) begin
        debug_7_36 = 1'b1;
      end else begin
        debug_7_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_295) begin
        debug_7_36 = 1'b1;
      end else begin
        debug_7_36 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_288 = (_zz_when_ArraySlice_l165_288 <= selectWriteFifo);
  assign when_ArraySlice_l166_288 = (_zz_when_ArraySlice_l166_288 <= _zz_when_ArraySlice_l166_288_1);
  assign _zz_when_ArraySlice_l112_288 = (wReg % _zz__zz_when_ArraySlice_l112_288);
  assign when_ArraySlice_l112_288 = (_zz_when_ArraySlice_l112_288 != 6'h0);
  assign when_ArraySlice_l113_288 = (7'h40 <= _zz_when_ArraySlice_l113_288);
  always @(*) begin
    if(when_ArraySlice_l112_288) begin
      if(when_ArraySlice_l113_288) begin
        _zz_when_ArraySlice_l173_288 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_288 = (_zz__zz_when_ArraySlice_l173_288 - _zz__zz_when_ArraySlice_l173_288_3);
      end
    end else begin
      if(when_ArraySlice_l118_288) begin
        _zz_when_ArraySlice_l173_288 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_288 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_288 = (_zz_when_ArraySlice_l118_288 <= wReg);
  assign when_ArraySlice_l173_288 = (_zz_when_ArraySlice_l173_288_1 <= _zz_when_ArraySlice_l173_288_2);
  assign when_ArraySlice_l165_289 = (_zz_when_ArraySlice_l165_289 <= selectWriteFifo);
  assign when_ArraySlice_l166_289 = (_zz_when_ArraySlice_l166_289 <= _zz_when_ArraySlice_l166_289_1);
  assign _zz_when_ArraySlice_l112_289 = (wReg % _zz__zz_when_ArraySlice_l112_289);
  assign when_ArraySlice_l112_289 = (_zz_when_ArraySlice_l112_289 != 6'h0);
  assign when_ArraySlice_l113_289 = (7'h40 <= _zz_when_ArraySlice_l113_289);
  always @(*) begin
    if(when_ArraySlice_l112_289) begin
      if(when_ArraySlice_l113_289) begin
        _zz_when_ArraySlice_l173_289 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_289 = (_zz__zz_when_ArraySlice_l173_289 - _zz__zz_when_ArraySlice_l173_289_3);
      end
    end else begin
      if(when_ArraySlice_l118_289) begin
        _zz_when_ArraySlice_l173_289 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_289 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_289 = (_zz_when_ArraySlice_l118_289 <= wReg);
  assign when_ArraySlice_l173_289 = (_zz_when_ArraySlice_l173_289_1 <= _zz_when_ArraySlice_l173_289_3);
  assign when_ArraySlice_l165_290 = (_zz_when_ArraySlice_l165_290 <= selectWriteFifo);
  assign when_ArraySlice_l166_290 = (_zz_when_ArraySlice_l166_290 <= _zz_when_ArraySlice_l166_290_1);
  assign _zz_when_ArraySlice_l112_290 = (wReg % _zz__zz_when_ArraySlice_l112_290);
  assign when_ArraySlice_l112_290 = (_zz_when_ArraySlice_l112_290 != 6'h0);
  assign when_ArraySlice_l113_290 = (7'h40 <= _zz_when_ArraySlice_l113_290);
  always @(*) begin
    if(when_ArraySlice_l112_290) begin
      if(when_ArraySlice_l113_290) begin
        _zz_when_ArraySlice_l173_290 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_290 = (_zz__zz_when_ArraySlice_l173_290 - _zz__zz_when_ArraySlice_l173_290_3);
      end
    end else begin
      if(when_ArraySlice_l118_290) begin
        _zz_when_ArraySlice_l173_290 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_290 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_290 = (_zz_when_ArraySlice_l118_290 <= wReg);
  assign when_ArraySlice_l173_290 = (_zz_when_ArraySlice_l173_290_1 <= _zz_when_ArraySlice_l173_290_3);
  assign when_ArraySlice_l165_291 = (_zz_when_ArraySlice_l165_291 <= selectWriteFifo);
  assign when_ArraySlice_l166_291 = (_zz_when_ArraySlice_l166_291 <= _zz_when_ArraySlice_l166_291_1);
  assign _zz_when_ArraySlice_l112_291 = (wReg % _zz__zz_when_ArraySlice_l112_291);
  assign when_ArraySlice_l112_291 = (_zz_when_ArraySlice_l112_291 != 6'h0);
  assign when_ArraySlice_l113_291 = (7'h40 <= _zz_when_ArraySlice_l113_291);
  always @(*) begin
    if(when_ArraySlice_l112_291) begin
      if(when_ArraySlice_l113_291) begin
        _zz_when_ArraySlice_l173_291 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_291 = (_zz__zz_when_ArraySlice_l173_291 - _zz__zz_when_ArraySlice_l173_291_3);
      end
    end else begin
      if(when_ArraySlice_l118_291) begin
        _zz_when_ArraySlice_l173_291 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_291 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_291 = (_zz_when_ArraySlice_l118_291 <= wReg);
  assign when_ArraySlice_l173_291 = (_zz_when_ArraySlice_l173_291_1 <= _zz_when_ArraySlice_l173_291_3);
  assign when_ArraySlice_l165_292 = (_zz_when_ArraySlice_l165_292 <= selectWriteFifo);
  assign when_ArraySlice_l166_292 = (_zz_when_ArraySlice_l166_292 <= _zz_when_ArraySlice_l166_292_1);
  assign _zz_when_ArraySlice_l112_292 = (wReg % _zz__zz_when_ArraySlice_l112_292);
  assign when_ArraySlice_l112_292 = (_zz_when_ArraySlice_l112_292 != 6'h0);
  assign when_ArraySlice_l113_292 = (7'h40 <= _zz_when_ArraySlice_l113_292);
  always @(*) begin
    if(when_ArraySlice_l112_292) begin
      if(when_ArraySlice_l113_292) begin
        _zz_when_ArraySlice_l173_292 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_292 = (_zz__zz_when_ArraySlice_l173_292 - _zz__zz_when_ArraySlice_l173_292_3);
      end
    end else begin
      if(when_ArraySlice_l118_292) begin
        _zz_when_ArraySlice_l173_292 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_292 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_292 = (_zz_when_ArraySlice_l118_292 <= wReg);
  assign when_ArraySlice_l173_292 = (_zz_when_ArraySlice_l173_292_1 <= _zz_when_ArraySlice_l173_292_3);
  assign when_ArraySlice_l165_293 = (_zz_when_ArraySlice_l165_293 <= selectWriteFifo);
  assign when_ArraySlice_l166_293 = (_zz_when_ArraySlice_l166_293 <= _zz_when_ArraySlice_l166_293_2);
  assign _zz_when_ArraySlice_l112_293 = (wReg % _zz__zz_when_ArraySlice_l112_293);
  assign when_ArraySlice_l112_293 = (_zz_when_ArraySlice_l112_293 != 6'h0);
  assign when_ArraySlice_l113_293 = (7'h40 <= _zz_when_ArraySlice_l113_293);
  always @(*) begin
    if(when_ArraySlice_l112_293) begin
      if(when_ArraySlice_l113_293) begin
        _zz_when_ArraySlice_l173_293 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_293 = (_zz__zz_when_ArraySlice_l173_293 - _zz__zz_when_ArraySlice_l173_293_3);
      end
    end else begin
      if(when_ArraySlice_l118_293) begin
        _zz_when_ArraySlice_l173_293 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_293 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_293 = (_zz_when_ArraySlice_l118_293 <= wReg);
  assign when_ArraySlice_l173_293 = (_zz_when_ArraySlice_l173_293_1 <= _zz_when_ArraySlice_l173_293_3);
  assign when_ArraySlice_l165_294 = (_zz_when_ArraySlice_l165_294 <= selectWriteFifo);
  assign when_ArraySlice_l166_294 = (_zz_when_ArraySlice_l166_294 <= _zz_when_ArraySlice_l166_294_2);
  assign _zz_when_ArraySlice_l112_294 = (wReg % _zz__zz_when_ArraySlice_l112_294);
  assign when_ArraySlice_l112_294 = (_zz_when_ArraySlice_l112_294 != 6'h0);
  assign when_ArraySlice_l113_294 = (7'h40 <= _zz_when_ArraySlice_l113_294);
  always @(*) begin
    if(when_ArraySlice_l112_294) begin
      if(when_ArraySlice_l113_294) begin
        _zz_when_ArraySlice_l173_294 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_294 = (_zz__zz_when_ArraySlice_l173_294 - _zz__zz_when_ArraySlice_l173_294_3);
      end
    end else begin
      if(when_ArraySlice_l118_294) begin
        _zz_when_ArraySlice_l173_294 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_294 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_294 = (_zz_when_ArraySlice_l118_294 <= wReg);
  assign when_ArraySlice_l173_294 = (_zz_when_ArraySlice_l173_294_1 <= _zz_when_ArraySlice_l173_294_3);
  assign when_ArraySlice_l165_295 = (_zz_when_ArraySlice_l165_295 <= selectWriteFifo);
  assign when_ArraySlice_l166_295 = (_zz_when_ArraySlice_l166_295 <= _zz_when_ArraySlice_l166_295_2);
  assign _zz_when_ArraySlice_l112_295 = (wReg % _zz__zz_when_ArraySlice_l112_295);
  assign when_ArraySlice_l112_295 = (_zz_when_ArraySlice_l112_295 != 6'h0);
  assign when_ArraySlice_l113_295 = (7'h40 <= _zz_when_ArraySlice_l113_295);
  always @(*) begin
    if(when_ArraySlice_l112_295) begin
      if(when_ArraySlice_l113_295) begin
        _zz_when_ArraySlice_l173_295 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_295 = (_zz__zz_when_ArraySlice_l173_295 - _zz__zz_when_ArraySlice_l173_295_3);
      end
    end else begin
      if(when_ArraySlice_l118_295) begin
        _zz_when_ArraySlice_l173_295 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_295 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_295 = (_zz_when_ArraySlice_l118_295 <= wReg);
  assign when_ArraySlice_l173_295 = (_zz_when_ArraySlice_l173_295_1 <= _zz_when_ArraySlice_l173_295_3);
  assign when_ArraySlice_l285_3 = (! ((((((_zz_when_ArraySlice_l285_3_1 && _zz_when_ArraySlice_l285_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l285_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l285_3_4 && _zz_when_ArraySlice_l285_3_5) && (debug_4_36 == _zz_when_ArraySlice_l285_3_6)) && (debug_5_36 == 1'b1)) && (debug_6_36 == 1'b1)) && (debug_7_36 == 1'b1))));
  assign when_ArraySlice_l288_3 = (wReg <= _zz_when_ArraySlice_l288_3_1);
  assign outputStreamArrayData_3_fire_10 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l292_3 = ((_zz_when_ArraySlice_l292_3_1 == 13'h0) && outputStreamArrayData_3_fire_10);
  assign outputStreamArrayData_3_fire_11 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l303_3 = ((handshakeTimes_3_value == _zz_when_ArraySlice_l303_3_1) && outputStreamArrayData_3_fire_11);
  assign _zz_when_ArraySlice_l94_35 = (hReg % _zz__zz_when_ArraySlice_l94_35);
  assign when_ArraySlice_l94_35 = (_zz_when_ArraySlice_l94_35 != 6'h0);
  assign when_ArraySlice_l95_35 = (7'h40 <= _zz_when_ArraySlice_l95_35);
  always @(*) begin
    if(when_ArraySlice_l94_35) begin
      if(when_ArraySlice_l95_35) begin
        _zz_when_ArraySlice_l304_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_3 = (_zz__zz_when_ArraySlice_l304_3_1 - _zz__zz_when_ArraySlice_l304_3_4);
      end
    end else begin
      if(when_ArraySlice_l99_35) begin
        _zz_when_ArraySlice_l304_3 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_3 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_35 = (_zz_when_ArraySlice_l99_35 <= hReg);
  assign when_ArraySlice_l304_3 = (_zz_when_ArraySlice_l304_3_1 < _zz_when_ArraySlice_l304_3_4);
  always @(*) begin
    debug_0_37 = 1'b0;
    if(when_ArraySlice_l165_296) begin
      if(when_ArraySlice_l166_296) begin
        debug_0_37 = 1'b1;
      end else begin
        debug_0_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_296) begin
        debug_0_37 = 1'b1;
      end else begin
        debug_0_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_37 = 1'b0;
    if(when_ArraySlice_l165_297) begin
      if(when_ArraySlice_l166_297) begin
        debug_1_37 = 1'b1;
      end else begin
        debug_1_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_297) begin
        debug_1_37 = 1'b1;
      end else begin
        debug_1_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_37 = 1'b0;
    if(when_ArraySlice_l165_298) begin
      if(when_ArraySlice_l166_298) begin
        debug_2_37 = 1'b1;
      end else begin
        debug_2_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_298) begin
        debug_2_37 = 1'b1;
      end else begin
        debug_2_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_37 = 1'b0;
    if(when_ArraySlice_l165_299) begin
      if(when_ArraySlice_l166_299) begin
        debug_3_37 = 1'b1;
      end else begin
        debug_3_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_299) begin
        debug_3_37 = 1'b1;
      end else begin
        debug_3_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_37 = 1'b0;
    if(when_ArraySlice_l165_300) begin
      if(when_ArraySlice_l166_300) begin
        debug_4_37 = 1'b1;
      end else begin
        debug_4_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_300) begin
        debug_4_37 = 1'b1;
      end else begin
        debug_4_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_37 = 1'b0;
    if(when_ArraySlice_l165_301) begin
      if(when_ArraySlice_l166_301) begin
        debug_5_37 = 1'b1;
      end else begin
        debug_5_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_301) begin
        debug_5_37 = 1'b1;
      end else begin
        debug_5_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_37 = 1'b0;
    if(when_ArraySlice_l165_302) begin
      if(when_ArraySlice_l166_302) begin
        debug_6_37 = 1'b1;
      end else begin
        debug_6_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_302) begin
        debug_6_37 = 1'b1;
      end else begin
        debug_6_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_37 = 1'b0;
    if(when_ArraySlice_l165_303) begin
      if(when_ArraySlice_l166_303) begin
        debug_7_37 = 1'b1;
      end else begin
        debug_7_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_303) begin
        debug_7_37 = 1'b1;
      end else begin
        debug_7_37 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_296 = (_zz_when_ArraySlice_l165_296 <= selectWriteFifo);
  assign when_ArraySlice_l166_296 = (_zz_when_ArraySlice_l166_296 <= _zz_when_ArraySlice_l166_296_1);
  assign _zz_when_ArraySlice_l112_296 = (wReg % _zz__zz_when_ArraySlice_l112_296);
  assign when_ArraySlice_l112_296 = (_zz_when_ArraySlice_l112_296 != 6'h0);
  assign when_ArraySlice_l113_296 = (7'h40 <= _zz_when_ArraySlice_l113_296);
  always @(*) begin
    if(when_ArraySlice_l112_296) begin
      if(when_ArraySlice_l113_296) begin
        _zz_when_ArraySlice_l173_296 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_296 = (_zz__zz_when_ArraySlice_l173_296 - _zz__zz_when_ArraySlice_l173_296_3);
      end
    end else begin
      if(when_ArraySlice_l118_296) begin
        _zz_when_ArraySlice_l173_296 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_296 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_296 = (_zz_when_ArraySlice_l118_296 <= wReg);
  assign when_ArraySlice_l173_296 = (_zz_when_ArraySlice_l173_296_1 <= _zz_when_ArraySlice_l173_296_2);
  assign when_ArraySlice_l165_297 = (_zz_when_ArraySlice_l165_297 <= selectWriteFifo);
  assign when_ArraySlice_l166_297 = (_zz_when_ArraySlice_l166_297 <= _zz_when_ArraySlice_l166_297_1);
  assign _zz_when_ArraySlice_l112_297 = (wReg % _zz__zz_when_ArraySlice_l112_297);
  assign when_ArraySlice_l112_297 = (_zz_when_ArraySlice_l112_297 != 6'h0);
  assign when_ArraySlice_l113_297 = (7'h40 <= _zz_when_ArraySlice_l113_297);
  always @(*) begin
    if(when_ArraySlice_l112_297) begin
      if(when_ArraySlice_l113_297) begin
        _zz_when_ArraySlice_l173_297 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_297 = (_zz__zz_when_ArraySlice_l173_297 - _zz__zz_when_ArraySlice_l173_297_3);
      end
    end else begin
      if(when_ArraySlice_l118_297) begin
        _zz_when_ArraySlice_l173_297 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_297 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_297 = (_zz_when_ArraySlice_l118_297 <= wReg);
  assign when_ArraySlice_l173_297 = (_zz_when_ArraySlice_l173_297_1 <= _zz_when_ArraySlice_l173_297_3);
  assign when_ArraySlice_l165_298 = (_zz_when_ArraySlice_l165_298 <= selectWriteFifo);
  assign when_ArraySlice_l166_298 = (_zz_when_ArraySlice_l166_298 <= _zz_when_ArraySlice_l166_298_1);
  assign _zz_when_ArraySlice_l112_298 = (wReg % _zz__zz_when_ArraySlice_l112_298);
  assign when_ArraySlice_l112_298 = (_zz_when_ArraySlice_l112_298 != 6'h0);
  assign when_ArraySlice_l113_298 = (7'h40 <= _zz_when_ArraySlice_l113_298);
  always @(*) begin
    if(when_ArraySlice_l112_298) begin
      if(when_ArraySlice_l113_298) begin
        _zz_when_ArraySlice_l173_298 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_298 = (_zz__zz_when_ArraySlice_l173_298 - _zz__zz_when_ArraySlice_l173_298_3);
      end
    end else begin
      if(when_ArraySlice_l118_298) begin
        _zz_when_ArraySlice_l173_298 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_298 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_298 = (_zz_when_ArraySlice_l118_298 <= wReg);
  assign when_ArraySlice_l173_298 = (_zz_when_ArraySlice_l173_298_1 <= _zz_when_ArraySlice_l173_298_3);
  assign when_ArraySlice_l165_299 = (_zz_when_ArraySlice_l165_299 <= selectWriteFifo);
  assign when_ArraySlice_l166_299 = (_zz_when_ArraySlice_l166_299 <= _zz_when_ArraySlice_l166_299_1);
  assign _zz_when_ArraySlice_l112_299 = (wReg % _zz__zz_when_ArraySlice_l112_299);
  assign when_ArraySlice_l112_299 = (_zz_when_ArraySlice_l112_299 != 6'h0);
  assign when_ArraySlice_l113_299 = (7'h40 <= _zz_when_ArraySlice_l113_299);
  always @(*) begin
    if(when_ArraySlice_l112_299) begin
      if(when_ArraySlice_l113_299) begin
        _zz_when_ArraySlice_l173_299 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_299 = (_zz__zz_when_ArraySlice_l173_299 - _zz__zz_when_ArraySlice_l173_299_3);
      end
    end else begin
      if(when_ArraySlice_l118_299) begin
        _zz_when_ArraySlice_l173_299 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_299 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_299 = (_zz_when_ArraySlice_l118_299 <= wReg);
  assign when_ArraySlice_l173_299 = (_zz_when_ArraySlice_l173_299_1 <= _zz_when_ArraySlice_l173_299_3);
  assign when_ArraySlice_l165_300 = (_zz_when_ArraySlice_l165_300 <= selectWriteFifo);
  assign when_ArraySlice_l166_300 = (_zz_when_ArraySlice_l166_300 <= _zz_when_ArraySlice_l166_300_1);
  assign _zz_when_ArraySlice_l112_300 = (wReg % _zz__zz_when_ArraySlice_l112_300);
  assign when_ArraySlice_l112_300 = (_zz_when_ArraySlice_l112_300 != 6'h0);
  assign when_ArraySlice_l113_300 = (7'h40 <= _zz_when_ArraySlice_l113_300);
  always @(*) begin
    if(when_ArraySlice_l112_300) begin
      if(when_ArraySlice_l113_300) begin
        _zz_when_ArraySlice_l173_300 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_300 = (_zz__zz_when_ArraySlice_l173_300 - _zz__zz_when_ArraySlice_l173_300_3);
      end
    end else begin
      if(when_ArraySlice_l118_300) begin
        _zz_when_ArraySlice_l173_300 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_300 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_300 = (_zz_when_ArraySlice_l118_300 <= wReg);
  assign when_ArraySlice_l173_300 = (_zz_when_ArraySlice_l173_300_1 <= _zz_when_ArraySlice_l173_300_3);
  assign when_ArraySlice_l165_301 = (_zz_when_ArraySlice_l165_301 <= selectWriteFifo);
  assign when_ArraySlice_l166_301 = (_zz_when_ArraySlice_l166_301 <= _zz_when_ArraySlice_l166_301_2);
  assign _zz_when_ArraySlice_l112_301 = (wReg % _zz__zz_when_ArraySlice_l112_301);
  assign when_ArraySlice_l112_301 = (_zz_when_ArraySlice_l112_301 != 6'h0);
  assign when_ArraySlice_l113_301 = (7'h40 <= _zz_when_ArraySlice_l113_301);
  always @(*) begin
    if(when_ArraySlice_l112_301) begin
      if(when_ArraySlice_l113_301) begin
        _zz_when_ArraySlice_l173_301 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_301 = (_zz__zz_when_ArraySlice_l173_301 - _zz__zz_when_ArraySlice_l173_301_3);
      end
    end else begin
      if(when_ArraySlice_l118_301) begin
        _zz_when_ArraySlice_l173_301 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_301 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_301 = (_zz_when_ArraySlice_l118_301 <= wReg);
  assign when_ArraySlice_l173_301 = (_zz_when_ArraySlice_l173_301_1 <= _zz_when_ArraySlice_l173_301_3);
  assign when_ArraySlice_l165_302 = (_zz_when_ArraySlice_l165_302 <= selectWriteFifo);
  assign when_ArraySlice_l166_302 = (_zz_when_ArraySlice_l166_302 <= _zz_when_ArraySlice_l166_302_2);
  assign _zz_when_ArraySlice_l112_302 = (wReg % _zz__zz_when_ArraySlice_l112_302);
  assign when_ArraySlice_l112_302 = (_zz_when_ArraySlice_l112_302 != 6'h0);
  assign when_ArraySlice_l113_302 = (7'h40 <= _zz_when_ArraySlice_l113_302);
  always @(*) begin
    if(when_ArraySlice_l112_302) begin
      if(when_ArraySlice_l113_302) begin
        _zz_when_ArraySlice_l173_302 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_302 = (_zz__zz_when_ArraySlice_l173_302 - _zz__zz_when_ArraySlice_l173_302_3);
      end
    end else begin
      if(when_ArraySlice_l118_302) begin
        _zz_when_ArraySlice_l173_302 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_302 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_302 = (_zz_when_ArraySlice_l118_302 <= wReg);
  assign when_ArraySlice_l173_302 = (_zz_when_ArraySlice_l173_302_1 <= _zz_when_ArraySlice_l173_302_3);
  assign when_ArraySlice_l165_303 = (_zz_when_ArraySlice_l165_303 <= selectWriteFifo);
  assign when_ArraySlice_l166_303 = (_zz_when_ArraySlice_l166_303 <= _zz_when_ArraySlice_l166_303_2);
  assign _zz_when_ArraySlice_l112_303 = (wReg % _zz__zz_when_ArraySlice_l112_303);
  assign when_ArraySlice_l112_303 = (_zz_when_ArraySlice_l112_303 != 6'h0);
  assign when_ArraySlice_l113_303 = (7'h40 <= _zz_when_ArraySlice_l113_303);
  always @(*) begin
    if(when_ArraySlice_l112_303) begin
      if(when_ArraySlice_l113_303) begin
        _zz_when_ArraySlice_l173_303 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_303 = (_zz__zz_when_ArraySlice_l173_303 - _zz__zz_when_ArraySlice_l173_303_3);
      end
    end else begin
      if(when_ArraySlice_l118_303) begin
        _zz_when_ArraySlice_l173_303 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_303 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_303 = (_zz_when_ArraySlice_l118_303 <= wReg);
  assign when_ArraySlice_l173_303 = (_zz_when_ArraySlice_l173_303_1 <= _zz_when_ArraySlice_l173_303_3);
  assign when_ArraySlice_l311_3 = (! ((((((_zz_when_ArraySlice_l311_3_1 && _zz_when_ArraySlice_l311_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l311_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l311_3_4 && _zz_when_ArraySlice_l311_3_5) && (debug_4_37 == _zz_when_ArraySlice_l311_3_6)) && (debug_5_37 == 1'b1)) && (debug_6_37 == 1'b1)) && (debug_7_37 == 1'b1))));
  assign outputStreamArrayData_3_fire_12 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l315_3 = ((_zz_when_ArraySlice_l315_3_1 == 13'h0) && outputStreamArrayData_3_fire_12);
  assign when_ArraySlice_l301_3 = (allowPadding_3 && (wReg <= _zz_when_ArraySlice_l301_3));
  assign outputStreamArrayData_3_fire_13 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l322_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l322_3_1);
  assign when_ArraySlice_l240_4 = (_zz_when_ArraySlice_l240_4 < wReg);
  assign when_ArraySlice_l241_4 = ((! holdReadOp_4) && (_zz_when_ArraySlice_l241_4 != 7'h0));
  assign _zz_outputStreamArrayData_4_valid_1 = (selectReadFifo_4 + _zz__zz_outputStreamArrayData_4_valid_1);
  assign _zz_15 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_4_valid_1);
  assign _zz_io_pop_ready_12 = outputStreamArrayData_4_ready;
  assign when_ArraySlice_l246_4 = (! holdReadOp_4);
  assign outputStreamArrayData_4_fire_7 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l247_4 = ((_zz_when_ArraySlice_l247_4_1 < _zz_when_ArraySlice_l247_4_3) && outputStreamArrayData_4_fire_7);
  assign when_ArraySlice_l248_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l248_4_1);
  assign when_ArraySlice_l251_4 = (_zz_when_ArraySlice_l251_4 == 13'h0);
  assign outputStreamArrayData_4_fire_8 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l256_4 = ((_zz_when_ArraySlice_l256_4_1 == _zz_when_ArraySlice_l256_4_4) && outputStreamArrayData_4_fire_8);
  assign when_ArraySlice_l257_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l257_4_1);
  assign _zz_when_ArraySlice_l94_36 = (hReg % _zz__zz_when_ArraySlice_l94_36);
  assign when_ArraySlice_l94_36 = (_zz_when_ArraySlice_l94_36 != 6'h0);
  assign when_ArraySlice_l95_36 = (7'h40 <= _zz_when_ArraySlice_l95_36);
  always @(*) begin
    if(when_ArraySlice_l94_36) begin
      if(when_ArraySlice_l95_36) begin
        _zz_when_ArraySlice_l259_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_4 = (_zz__zz_when_ArraySlice_l259_4 - _zz__zz_when_ArraySlice_l259_4_3);
      end
    end else begin
      if(when_ArraySlice_l99_36) begin
        _zz_when_ArraySlice_l259_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_4 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_36 = (_zz_when_ArraySlice_l99_36 <= hReg);
  assign when_ArraySlice_l259_4 = (_zz_when_ArraySlice_l259_4_1 < _zz_when_ArraySlice_l259_4_4);
  always @(*) begin
    debug_0_38 = 1'b0;
    if(when_ArraySlice_l165_304) begin
      if(when_ArraySlice_l166_304) begin
        debug_0_38 = 1'b1;
      end else begin
        debug_0_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_304) begin
        debug_0_38 = 1'b1;
      end else begin
        debug_0_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_38 = 1'b0;
    if(when_ArraySlice_l165_305) begin
      if(when_ArraySlice_l166_305) begin
        debug_1_38 = 1'b1;
      end else begin
        debug_1_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_305) begin
        debug_1_38 = 1'b1;
      end else begin
        debug_1_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_38 = 1'b0;
    if(when_ArraySlice_l165_306) begin
      if(when_ArraySlice_l166_306) begin
        debug_2_38 = 1'b1;
      end else begin
        debug_2_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_306) begin
        debug_2_38 = 1'b1;
      end else begin
        debug_2_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_38 = 1'b0;
    if(when_ArraySlice_l165_307) begin
      if(when_ArraySlice_l166_307) begin
        debug_3_38 = 1'b1;
      end else begin
        debug_3_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_307) begin
        debug_3_38 = 1'b1;
      end else begin
        debug_3_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_38 = 1'b0;
    if(when_ArraySlice_l165_308) begin
      if(when_ArraySlice_l166_308) begin
        debug_4_38 = 1'b1;
      end else begin
        debug_4_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_308) begin
        debug_4_38 = 1'b1;
      end else begin
        debug_4_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_38 = 1'b0;
    if(when_ArraySlice_l165_309) begin
      if(when_ArraySlice_l166_309) begin
        debug_5_38 = 1'b1;
      end else begin
        debug_5_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_309) begin
        debug_5_38 = 1'b1;
      end else begin
        debug_5_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_38 = 1'b0;
    if(when_ArraySlice_l165_310) begin
      if(when_ArraySlice_l166_310) begin
        debug_6_38 = 1'b1;
      end else begin
        debug_6_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_310) begin
        debug_6_38 = 1'b1;
      end else begin
        debug_6_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_38 = 1'b0;
    if(when_ArraySlice_l165_311) begin
      if(when_ArraySlice_l166_311) begin
        debug_7_38 = 1'b1;
      end else begin
        debug_7_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_311) begin
        debug_7_38 = 1'b1;
      end else begin
        debug_7_38 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_304 = (_zz_when_ArraySlice_l165_304 <= selectWriteFifo);
  assign when_ArraySlice_l166_304 = (_zz_when_ArraySlice_l166_304 <= _zz_when_ArraySlice_l166_304_1);
  assign _zz_when_ArraySlice_l112_304 = (wReg % _zz__zz_when_ArraySlice_l112_304);
  assign when_ArraySlice_l112_304 = (_zz_when_ArraySlice_l112_304 != 6'h0);
  assign when_ArraySlice_l113_304 = (7'h40 <= _zz_when_ArraySlice_l113_304);
  always @(*) begin
    if(when_ArraySlice_l112_304) begin
      if(when_ArraySlice_l113_304) begin
        _zz_when_ArraySlice_l173_304 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_304 = (_zz__zz_when_ArraySlice_l173_304 - _zz__zz_when_ArraySlice_l173_304_3);
      end
    end else begin
      if(when_ArraySlice_l118_304) begin
        _zz_when_ArraySlice_l173_304 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_304 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_304 = (_zz_when_ArraySlice_l118_304 <= wReg);
  assign when_ArraySlice_l173_304 = (_zz_when_ArraySlice_l173_304_1 <= _zz_when_ArraySlice_l173_304_2);
  assign when_ArraySlice_l165_305 = (_zz_when_ArraySlice_l165_305 <= selectWriteFifo);
  assign when_ArraySlice_l166_305 = (_zz_when_ArraySlice_l166_305 <= _zz_when_ArraySlice_l166_305_1);
  assign _zz_when_ArraySlice_l112_305 = (wReg % _zz__zz_when_ArraySlice_l112_305);
  assign when_ArraySlice_l112_305 = (_zz_when_ArraySlice_l112_305 != 6'h0);
  assign when_ArraySlice_l113_305 = (7'h40 <= _zz_when_ArraySlice_l113_305);
  always @(*) begin
    if(when_ArraySlice_l112_305) begin
      if(when_ArraySlice_l113_305) begin
        _zz_when_ArraySlice_l173_305 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_305 = (_zz__zz_when_ArraySlice_l173_305 - _zz__zz_when_ArraySlice_l173_305_3);
      end
    end else begin
      if(when_ArraySlice_l118_305) begin
        _zz_when_ArraySlice_l173_305 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_305 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_305 = (_zz_when_ArraySlice_l118_305 <= wReg);
  assign when_ArraySlice_l173_305 = (_zz_when_ArraySlice_l173_305_1 <= _zz_when_ArraySlice_l173_305_3);
  assign when_ArraySlice_l165_306 = (_zz_when_ArraySlice_l165_306 <= selectWriteFifo);
  assign when_ArraySlice_l166_306 = (_zz_when_ArraySlice_l166_306 <= _zz_when_ArraySlice_l166_306_1);
  assign _zz_when_ArraySlice_l112_306 = (wReg % _zz__zz_when_ArraySlice_l112_306);
  assign when_ArraySlice_l112_306 = (_zz_when_ArraySlice_l112_306 != 6'h0);
  assign when_ArraySlice_l113_306 = (7'h40 <= _zz_when_ArraySlice_l113_306);
  always @(*) begin
    if(when_ArraySlice_l112_306) begin
      if(when_ArraySlice_l113_306) begin
        _zz_when_ArraySlice_l173_306 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_306 = (_zz__zz_when_ArraySlice_l173_306 - _zz__zz_when_ArraySlice_l173_306_3);
      end
    end else begin
      if(when_ArraySlice_l118_306) begin
        _zz_when_ArraySlice_l173_306 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_306 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_306 = (_zz_when_ArraySlice_l118_306 <= wReg);
  assign when_ArraySlice_l173_306 = (_zz_when_ArraySlice_l173_306_1 <= _zz_when_ArraySlice_l173_306_3);
  assign when_ArraySlice_l165_307 = (_zz_when_ArraySlice_l165_307 <= selectWriteFifo);
  assign when_ArraySlice_l166_307 = (_zz_when_ArraySlice_l166_307 <= _zz_when_ArraySlice_l166_307_1);
  assign _zz_when_ArraySlice_l112_307 = (wReg % _zz__zz_when_ArraySlice_l112_307);
  assign when_ArraySlice_l112_307 = (_zz_when_ArraySlice_l112_307 != 6'h0);
  assign when_ArraySlice_l113_307 = (7'h40 <= _zz_when_ArraySlice_l113_307);
  always @(*) begin
    if(when_ArraySlice_l112_307) begin
      if(when_ArraySlice_l113_307) begin
        _zz_when_ArraySlice_l173_307 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_307 = (_zz__zz_when_ArraySlice_l173_307 - _zz__zz_when_ArraySlice_l173_307_3);
      end
    end else begin
      if(when_ArraySlice_l118_307) begin
        _zz_when_ArraySlice_l173_307 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_307 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_307 = (_zz_when_ArraySlice_l118_307 <= wReg);
  assign when_ArraySlice_l173_307 = (_zz_when_ArraySlice_l173_307_1 <= _zz_when_ArraySlice_l173_307_3);
  assign when_ArraySlice_l165_308 = (_zz_when_ArraySlice_l165_308 <= selectWriteFifo);
  assign when_ArraySlice_l166_308 = (_zz_when_ArraySlice_l166_308 <= _zz_when_ArraySlice_l166_308_1);
  assign _zz_when_ArraySlice_l112_308 = (wReg % _zz__zz_when_ArraySlice_l112_308);
  assign when_ArraySlice_l112_308 = (_zz_when_ArraySlice_l112_308 != 6'h0);
  assign when_ArraySlice_l113_308 = (7'h40 <= _zz_when_ArraySlice_l113_308);
  always @(*) begin
    if(when_ArraySlice_l112_308) begin
      if(when_ArraySlice_l113_308) begin
        _zz_when_ArraySlice_l173_308 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_308 = (_zz__zz_when_ArraySlice_l173_308 - _zz__zz_when_ArraySlice_l173_308_3);
      end
    end else begin
      if(when_ArraySlice_l118_308) begin
        _zz_when_ArraySlice_l173_308 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_308 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_308 = (_zz_when_ArraySlice_l118_308 <= wReg);
  assign when_ArraySlice_l173_308 = (_zz_when_ArraySlice_l173_308_1 <= _zz_when_ArraySlice_l173_308_3);
  assign when_ArraySlice_l165_309 = (_zz_when_ArraySlice_l165_309 <= selectWriteFifo);
  assign when_ArraySlice_l166_309 = (_zz_when_ArraySlice_l166_309 <= _zz_when_ArraySlice_l166_309_2);
  assign _zz_when_ArraySlice_l112_309 = (wReg % _zz__zz_when_ArraySlice_l112_309);
  assign when_ArraySlice_l112_309 = (_zz_when_ArraySlice_l112_309 != 6'h0);
  assign when_ArraySlice_l113_309 = (7'h40 <= _zz_when_ArraySlice_l113_309);
  always @(*) begin
    if(when_ArraySlice_l112_309) begin
      if(when_ArraySlice_l113_309) begin
        _zz_when_ArraySlice_l173_309 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_309 = (_zz__zz_when_ArraySlice_l173_309 - _zz__zz_when_ArraySlice_l173_309_3);
      end
    end else begin
      if(when_ArraySlice_l118_309) begin
        _zz_when_ArraySlice_l173_309 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_309 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_309 = (_zz_when_ArraySlice_l118_309 <= wReg);
  assign when_ArraySlice_l173_309 = (_zz_when_ArraySlice_l173_309_1 <= _zz_when_ArraySlice_l173_309_3);
  assign when_ArraySlice_l165_310 = (_zz_when_ArraySlice_l165_310 <= selectWriteFifo);
  assign when_ArraySlice_l166_310 = (_zz_when_ArraySlice_l166_310 <= _zz_when_ArraySlice_l166_310_2);
  assign _zz_when_ArraySlice_l112_310 = (wReg % _zz__zz_when_ArraySlice_l112_310);
  assign when_ArraySlice_l112_310 = (_zz_when_ArraySlice_l112_310 != 6'h0);
  assign when_ArraySlice_l113_310 = (7'h40 <= _zz_when_ArraySlice_l113_310);
  always @(*) begin
    if(when_ArraySlice_l112_310) begin
      if(when_ArraySlice_l113_310) begin
        _zz_when_ArraySlice_l173_310 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_310 = (_zz__zz_when_ArraySlice_l173_310 - _zz__zz_when_ArraySlice_l173_310_3);
      end
    end else begin
      if(when_ArraySlice_l118_310) begin
        _zz_when_ArraySlice_l173_310 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_310 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_310 = (_zz_when_ArraySlice_l118_310 <= wReg);
  assign when_ArraySlice_l173_310 = (_zz_when_ArraySlice_l173_310_1 <= _zz_when_ArraySlice_l173_310_3);
  assign when_ArraySlice_l165_311 = (_zz_when_ArraySlice_l165_311 <= selectWriteFifo);
  assign when_ArraySlice_l166_311 = (_zz_when_ArraySlice_l166_311 <= _zz_when_ArraySlice_l166_311_2);
  assign _zz_when_ArraySlice_l112_311 = (wReg % _zz__zz_when_ArraySlice_l112_311);
  assign when_ArraySlice_l112_311 = (_zz_when_ArraySlice_l112_311 != 6'h0);
  assign when_ArraySlice_l113_311 = (7'h40 <= _zz_when_ArraySlice_l113_311);
  always @(*) begin
    if(when_ArraySlice_l112_311) begin
      if(when_ArraySlice_l113_311) begin
        _zz_when_ArraySlice_l173_311 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_311 = (_zz__zz_when_ArraySlice_l173_311 - _zz__zz_when_ArraySlice_l173_311_3);
      end
    end else begin
      if(when_ArraySlice_l118_311) begin
        _zz_when_ArraySlice_l173_311 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_311 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_311 = (_zz_when_ArraySlice_l118_311 <= wReg);
  assign when_ArraySlice_l173_311 = (_zz_when_ArraySlice_l173_311_1 <= _zz_when_ArraySlice_l173_311_3);
  assign when_ArraySlice_l265_4 = (! ((((((_zz_when_ArraySlice_l265_4_1 && _zz_when_ArraySlice_l265_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l265_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l265_4_4 && _zz_when_ArraySlice_l265_4_5) && (debug_4_38 == _zz_when_ArraySlice_l265_4_6)) && (debug_5_38 == 1'b1)) && (debug_6_38 == 1'b1)) && (debug_7_38 == 1'b1))));
  assign when_ArraySlice_l268_4 = (wReg <= _zz_when_ArraySlice_l268_4_1);
  assign when_ArraySlice_l272_4 = (_zz_when_ArraySlice_l272_4 == 13'h0);
  assign when_ArraySlice_l276_4 = (_zz_when_ArraySlice_l276_4 == 7'h0);
  assign outputStreamArrayData_4_fire_9 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l277_4 = ((handshakeTimes_4_value == _zz_when_ArraySlice_l277_4_1) && outputStreamArrayData_4_fire_9);
  assign _zz_when_ArraySlice_l94_37 = (hReg % _zz__zz_when_ArraySlice_l94_37);
  assign when_ArraySlice_l94_37 = (_zz_when_ArraySlice_l94_37 != 6'h0);
  assign when_ArraySlice_l95_37 = (7'h40 <= _zz_when_ArraySlice_l95_37);
  always @(*) begin
    if(when_ArraySlice_l94_37) begin
      if(when_ArraySlice_l95_37) begin
        _zz_when_ArraySlice_l279_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_4 = (_zz__zz_when_ArraySlice_l279_4 - _zz__zz_when_ArraySlice_l279_4_3);
      end
    end else begin
      if(when_ArraySlice_l99_37) begin
        _zz_when_ArraySlice_l279_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_4 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_37 = (_zz_when_ArraySlice_l99_37 <= hReg);
  assign when_ArraySlice_l279_4 = (_zz_when_ArraySlice_l279_4_1 < _zz_when_ArraySlice_l279_4_4);
  always @(*) begin
    debug_0_39 = 1'b0;
    if(when_ArraySlice_l165_312) begin
      if(when_ArraySlice_l166_312) begin
        debug_0_39 = 1'b1;
      end else begin
        debug_0_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_312) begin
        debug_0_39 = 1'b1;
      end else begin
        debug_0_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_39 = 1'b0;
    if(when_ArraySlice_l165_313) begin
      if(when_ArraySlice_l166_313) begin
        debug_1_39 = 1'b1;
      end else begin
        debug_1_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_313) begin
        debug_1_39 = 1'b1;
      end else begin
        debug_1_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_39 = 1'b0;
    if(when_ArraySlice_l165_314) begin
      if(when_ArraySlice_l166_314) begin
        debug_2_39 = 1'b1;
      end else begin
        debug_2_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_314) begin
        debug_2_39 = 1'b1;
      end else begin
        debug_2_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_39 = 1'b0;
    if(when_ArraySlice_l165_315) begin
      if(when_ArraySlice_l166_315) begin
        debug_3_39 = 1'b1;
      end else begin
        debug_3_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_315) begin
        debug_3_39 = 1'b1;
      end else begin
        debug_3_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_39 = 1'b0;
    if(when_ArraySlice_l165_316) begin
      if(when_ArraySlice_l166_316) begin
        debug_4_39 = 1'b1;
      end else begin
        debug_4_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_316) begin
        debug_4_39 = 1'b1;
      end else begin
        debug_4_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_39 = 1'b0;
    if(when_ArraySlice_l165_317) begin
      if(when_ArraySlice_l166_317) begin
        debug_5_39 = 1'b1;
      end else begin
        debug_5_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_317) begin
        debug_5_39 = 1'b1;
      end else begin
        debug_5_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_39 = 1'b0;
    if(when_ArraySlice_l165_318) begin
      if(when_ArraySlice_l166_318) begin
        debug_6_39 = 1'b1;
      end else begin
        debug_6_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_318) begin
        debug_6_39 = 1'b1;
      end else begin
        debug_6_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_39 = 1'b0;
    if(when_ArraySlice_l165_319) begin
      if(when_ArraySlice_l166_319) begin
        debug_7_39 = 1'b1;
      end else begin
        debug_7_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_319) begin
        debug_7_39 = 1'b1;
      end else begin
        debug_7_39 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_312 = (_zz_when_ArraySlice_l165_312 <= selectWriteFifo);
  assign when_ArraySlice_l166_312 = (_zz_when_ArraySlice_l166_312 <= _zz_when_ArraySlice_l166_312_1);
  assign _zz_when_ArraySlice_l112_312 = (wReg % _zz__zz_when_ArraySlice_l112_312);
  assign when_ArraySlice_l112_312 = (_zz_when_ArraySlice_l112_312 != 6'h0);
  assign when_ArraySlice_l113_312 = (7'h40 <= _zz_when_ArraySlice_l113_312);
  always @(*) begin
    if(when_ArraySlice_l112_312) begin
      if(when_ArraySlice_l113_312) begin
        _zz_when_ArraySlice_l173_312 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_312 = (_zz__zz_when_ArraySlice_l173_312 - _zz__zz_when_ArraySlice_l173_312_3);
      end
    end else begin
      if(when_ArraySlice_l118_312) begin
        _zz_when_ArraySlice_l173_312 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_312 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_312 = (_zz_when_ArraySlice_l118_312 <= wReg);
  assign when_ArraySlice_l173_312 = (_zz_when_ArraySlice_l173_312_1 <= _zz_when_ArraySlice_l173_312_2);
  assign when_ArraySlice_l165_313 = (_zz_when_ArraySlice_l165_313 <= selectWriteFifo);
  assign when_ArraySlice_l166_313 = (_zz_when_ArraySlice_l166_313 <= _zz_when_ArraySlice_l166_313_1);
  assign _zz_when_ArraySlice_l112_313 = (wReg % _zz__zz_when_ArraySlice_l112_313);
  assign when_ArraySlice_l112_313 = (_zz_when_ArraySlice_l112_313 != 6'h0);
  assign when_ArraySlice_l113_313 = (7'h40 <= _zz_when_ArraySlice_l113_313);
  always @(*) begin
    if(when_ArraySlice_l112_313) begin
      if(when_ArraySlice_l113_313) begin
        _zz_when_ArraySlice_l173_313 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_313 = (_zz__zz_when_ArraySlice_l173_313 - _zz__zz_when_ArraySlice_l173_313_3);
      end
    end else begin
      if(when_ArraySlice_l118_313) begin
        _zz_when_ArraySlice_l173_313 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_313 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_313 = (_zz_when_ArraySlice_l118_313 <= wReg);
  assign when_ArraySlice_l173_313 = (_zz_when_ArraySlice_l173_313_1 <= _zz_when_ArraySlice_l173_313_3);
  assign when_ArraySlice_l165_314 = (_zz_when_ArraySlice_l165_314 <= selectWriteFifo);
  assign when_ArraySlice_l166_314 = (_zz_when_ArraySlice_l166_314 <= _zz_when_ArraySlice_l166_314_1);
  assign _zz_when_ArraySlice_l112_314 = (wReg % _zz__zz_when_ArraySlice_l112_314);
  assign when_ArraySlice_l112_314 = (_zz_when_ArraySlice_l112_314 != 6'h0);
  assign when_ArraySlice_l113_314 = (7'h40 <= _zz_when_ArraySlice_l113_314);
  always @(*) begin
    if(when_ArraySlice_l112_314) begin
      if(when_ArraySlice_l113_314) begin
        _zz_when_ArraySlice_l173_314 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_314 = (_zz__zz_when_ArraySlice_l173_314 - _zz__zz_when_ArraySlice_l173_314_3);
      end
    end else begin
      if(when_ArraySlice_l118_314) begin
        _zz_when_ArraySlice_l173_314 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_314 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_314 = (_zz_when_ArraySlice_l118_314 <= wReg);
  assign when_ArraySlice_l173_314 = (_zz_when_ArraySlice_l173_314_1 <= _zz_when_ArraySlice_l173_314_3);
  assign when_ArraySlice_l165_315 = (_zz_when_ArraySlice_l165_315 <= selectWriteFifo);
  assign when_ArraySlice_l166_315 = (_zz_when_ArraySlice_l166_315 <= _zz_when_ArraySlice_l166_315_1);
  assign _zz_when_ArraySlice_l112_315 = (wReg % _zz__zz_when_ArraySlice_l112_315);
  assign when_ArraySlice_l112_315 = (_zz_when_ArraySlice_l112_315 != 6'h0);
  assign when_ArraySlice_l113_315 = (7'h40 <= _zz_when_ArraySlice_l113_315);
  always @(*) begin
    if(when_ArraySlice_l112_315) begin
      if(when_ArraySlice_l113_315) begin
        _zz_when_ArraySlice_l173_315 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_315 = (_zz__zz_when_ArraySlice_l173_315 - _zz__zz_when_ArraySlice_l173_315_3);
      end
    end else begin
      if(when_ArraySlice_l118_315) begin
        _zz_when_ArraySlice_l173_315 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_315 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_315 = (_zz_when_ArraySlice_l118_315 <= wReg);
  assign when_ArraySlice_l173_315 = (_zz_when_ArraySlice_l173_315_1 <= _zz_when_ArraySlice_l173_315_3);
  assign when_ArraySlice_l165_316 = (_zz_when_ArraySlice_l165_316 <= selectWriteFifo);
  assign when_ArraySlice_l166_316 = (_zz_when_ArraySlice_l166_316 <= _zz_when_ArraySlice_l166_316_1);
  assign _zz_when_ArraySlice_l112_316 = (wReg % _zz__zz_when_ArraySlice_l112_316);
  assign when_ArraySlice_l112_316 = (_zz_when_ArraySlice_l112_316 != 6'h0);
  assign when_ArraySlice_l113_316 = (7'h40 <= _zz_when_ArraySlice_l113_316);
  always @(*) begin
    if(when_ArraySlice_l112_316) begin
      if(when_ArraySlice_l113_316) begin
        _zz_when_ArraySlice_l173_316 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_316 = (_zz__zz_when_ArraySlice_l173_316 - _zz__zz_when_ArraySlice_l173_316_3);
      end
    end else begin
      if(when_ArraySlice_l118_316) begin
        _zz_when_ArraySlice_l173_316 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_316 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_316 = (_zz_when_ArraySlice_l118_316 <= wReg);
  assign when_ArraySlice_l173_316 = (_zz_when_ArraySlice_l173_316_1 <= _zz_when_ArraySlice_l173_316_3);
  assign when_ArraySlice_l165_317 = (_zz_when_ArraySlice_l165_317 <= selectWriteFifo);
  assign when_ArraySlice_l166_317 = (_zz_when_ArraySlice_l166_317 <= _zz_when_ArraySlice_l166_317_2);
  assign _zz_when_ArraySlice_l112_317 = (wReg % _zz__zz_when_ArraySlice_l112_317);
  assign when_ArraySlice_l112_317 = (_zz_when_ArraySlice_l112_317 != 6'h0);
  assign when_ArraySlice_l113_317 = (7'h40 <= _zz_when_ArraySlice_l113_317);
  always @(*) begin
    if(when_ArraySlice_l112_317) begin
      if(when_ArraySlice_l113_317) begin
        _zz_when_ArraySlice_l173_317 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_317 = (_zz__zz_when_ArraySlice_l173_317 - _zz__zz_when_ArraySlice_l173_317_3);
      end
    end else begin
      if(when_ArraySlice_l118_317) begin
        _zz_when_ArraySlice_l173_317 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_317 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_317 = (_zz_when_ArraySlice_l118_317 <= wReg);
  assign when_ArraySlice_l173_317 = (_zz_when_ArraySlice_l173_317_1 <= _zz_when_ArraySlice_l173_317_3);
  assign when_ArraySlice_l165_318 = (_zz_when_ArraySlice_l165_318 <= selectWriteFifo);
  assign when_ArraySlice_l166_318 = (_zz_when_ArraySlice_l166_318 <= _zz_when_ArraySlice_l166_318_2);
  assign _zz_when_ArraySlice_l112_318 = (wReg % _zz__zz_when_ArraySlice_l112_318);
  assign when_ArraySlice_l112_318 = (_zz_when_ArraySlice_l112_318 != 6'h0);
  assign when_ArraySlice_l113_318 = (7'h40 <= _zz_when_ArraySlice_l113_318);
  always @(*) begin
    if(when_ArraySlice_l112_318) begin
      if(when_ArraySlice_l113_318) begin
        _zz_when_ArraySlice_l173_318 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_318 = (_zz__zz_when_ArraySlice_l173_318 - _zz__zz_when_ArraySlice_l173_318_3);
      end
    end else begin
      if(when_ArraySlice_l118_318) begin
        _zz_when_ArraySlice_l173_318 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_318 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_318 = (_zz_when_ArraySlice_l118_318 <= wReg);
  assign when_ArraySlice_l173_318 = (_zz_when_ArraySlice_l173_318_1 <= _zz_when_ArraySlice_l173_318_3);
  assign when_ArraySlice_l165_319 = (_zz_when_ArraySlice_l165_319 <= selectWriteFifo);
  assign when_ArraySlice_l166_319 = (_zz_when_ArraySlice_l166_319 <= _zz_when_ArraySlice_l166_319_2);
  assign _zz_when_ArraySlice_l112_319 = (wReg % _zz__zz_when_ArraySlice_l112_319);
  assign when_ArraySlice_l112_319 = (_zz_when_ArraySlice_l112_319 != 6'h0);
  assign when_ArraySlice_l113_319 = (7'h40 <= _zz_when_ArraySlice_l113_319);
  always @(*) begin
    if(when_ArraySlice_l112_319) begin
      if(when_ArraySlice_l113_319) begin
        _zz_when_ArraySlice_l173_319 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_319 = (_zz__zz_when_ArraySlice_l173_319 - _zz__zz_when_ArraySlice_l173_319_3);
      end
    end else begin
      if(when_ArraySlice_l118_319) begin
        _zz_when_ArraySlice_l173_319 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_319 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_319 = (_zz_when_ArraySlice_l118_319 <= wReg);
  assign when_ArraySlice_l173_319 = (_zz_when_ArraySlice_l173_319_1 <= _zz_when_ArraySlice_l173_319_3);
  assign when_ArraySlice_l285_4 = (! ((((((_zz_when_ArraySlice_l285_4_1 && _zz_when_ArraySlice_l285_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l285_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l285_4_4 && _zz_when_ArraySlice_l285_4_5) && (debug_4_39 == _zz_when_ArraySlice_l285_4_6)) && (debug_5_39 == 1'b1)) && (debug_6_39 == 1'b1)) && (debug_7_39 == 1'b1))));
  assign when_ArraySlice_l288_4 = (wReg <= _zz_when_ArraySlice_l288_4_1);
  assign outputStreamArrayData_4_fire_10 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l292_4 = ((_zz_when_ArraySlice_l292_4 == 13'h0) && outputStreamArrayData_4_fire_10);
  assign outputStreamArrayData_4_fire_11 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l303_4 = ((handshakeTimes_4_value == _zz_when_ArraySlice_l303_4_1) && outputStreamArrayData_4_fire_11);
  assign _zz_when_ArraySlice_l94_38 = (hReg % _zz__zz_when_ArraySlice_l94_38);
  assign when_ArraySlice_l94_38 = (_zz_when_ArraySlice_l94_38 != 6'h0);
  assign when_ArraySlice_l95_38 = (7'h40 <= _zz_when_ArraySlice_l95_38);
  always @(*) begin
    if(when_ArraySlice_l94_38) begin
      if(when_ArraySlice_l95_38) begin
        _zz_when_ArraySlice_l304_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_4 = (_zz__zz_when_ArraySlice_l304_4 - _zz__zz_when_ArraySlice_l304_4_3);
      end
    end else begin
      if(when_ArraySlice_l99_38) begin
        _zz_when_ArraySlice_l304_4 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_4 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_38 = (_zz_when_ArraySlice_l99_38 <= hReg);
  assign when_ArraySlice_l304_4 = (_zz_when_ArraySlice_l304_4_1 < _zz_when_ArraySlice_l304_4_4);
  always @(*) begin
    debug_0_40 = 1'b0;
    if(when_ArraySlice_l165_320) begin
      if(when_ArraySlice_l166_320) begin
        debug_0_40 = 1'b1;
      end else begin
        debug_0_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_320) begin
        debug_0_40 = 1'b1;
      end else begin
        debug_0_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_40 = 1'b0;
    if(when_ArraySlice_l165_321) begin
      if(when_ArraySlice_l166_321) begin
        debug_1_40 = 1'b1;
      end else begin
        debug_1_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_321) begin
        debug_1_40 = 1'b1;
      end else begin
        debug_1_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_40 = 1'b0;
    if(when_ArraySlice_l165_322) begin
      if(when_ArraySlice_l166_322) begin
        debug_2_40 = 1'b1;
      end else begin
        debug_2_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_322) begin
        debug_2_40 = 1'b1;
      end else begin
        debug_2_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_40 = 1'b0;
    if(when_ArraySlice_l165_323) begin
      if(when_ArraySlice_l166_323) begin
        debug_3_40 = 1'b1;
      end else begin
        debug_3_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_323) begin
        debug_3_40 = 1'b1;
      end else begin
        debug_3_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_40 = 1'b0;
    if(when_ArraySlice_l165_324) begin
      if(when_ArraySlice_l166_324) begin
        debug_4_40 = 1'b1;
      end else begin
        debug_4_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_324) begin
        debug_4_40 = 1'b1;
      end else begin
        debug_4_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_40 = 1'b0;
    if(when_ArraySlice_l165_325) begin
      if(when_ArraySlice_l166_325) begin
        debug_5_40 = 1'b1;
      end else begin
        debug_5_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_325) begin
        debug_5_40 = 1'b1;
      end else begin
        debug_5_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_40 = 1'b0;
    if(when_ArraySlice_l165_326) begin
      if(when_ArraySlice_l166_326) begin
        debug_6_40 = 1'b1;
      end else begin
        debug_6_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_326) begin
        debug_6_40 = 1'b1;
      end else begin
        debug_6_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_40 = 1'b0;
    if(when_ArraySlice_l165_327) begin
      if(when_ArraySlice_l166_327) begin
        debug_7_40 = 1'b1;
      end else begin
        debug_7_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_327) begin
        debug_7_40 = 1'b1;
      end else begin
        debug_7_40 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_320 = (_zz_when_ArraySlice_l165_320 <= selectWriteFifo);
  assign when_ArraySlice_l166_320 = (_zz_when_ArraySlice_l166_320 <= _zz_when_ArraySlice_l166_320_1);
  assign _zz_when_ArraySlice_l112_320 = (wReg % _zz__zz_when_ArraySlice_l112_320);
  assign when_ArraySlice_l112_320 = (_zz_when_ArraySlice_l112_320 != 6'h0);
  assign when_ArraySlice_l113_320 = (7'h40 <= _zz_when_ArraySlice_l113_320);
  always @(*) begin
    if(when_ArraySlice_l112_320) begin
      if(when_ArraySlice_l113_320) begin
        _zz_when_ArraySlice_l173_320 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_320 = (_zz__zz_when_ArraySlice_l173_320 - _zz__zz_when_ArraySlice_l173_320_3);
      end
    end else begin
      if(when_ArraySlice_l118_320) begin
        _zz_when_ArraySlice_l173_320 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_320 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_320 = (_zz_when_ArraySlice_l118_320 <= wReg);
  assign when_ArraySlice_l173_320 = (_zz_when_ArraySlice_l173_320_1 <= _zz_when_ArraySlice_l173_320_2);
  assign when_ArraySlice_l165_321 = (_zz_when_ArraySlice_l165_321 <= selectWriteFifo);
  assign when_ArraySlice_l166_321 = (_zz_when_ArraySlice_l166_321 <= _zz_when_ArraySlice_l166_321_1);
  assign _zz_when_ArraySlice_l112_321 = (wReg % _zz__zz_when_ArraySlice_l112_321);
  assign when_ArraySlice_l112_321 = (_zz_when_ArraySlice_l112_321 != 6'h0);
  assign when_ArraySlice_l113_321 = (7'h40 <= _zz_when_ArraySlice_l113_321);
  always @(*) begin
    if(when_ArraySlice_l112_321) begin
      if(when_ArraySlice_l113_321) begin
        _zz_when_ArraySlice_l173_321 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_321 = (_zz__zz_when_ArraySlice_l173_321 - _zz__zz_when_ArraySlice_l173_321_3);
      end
    end else begin
      if(when_ArraySlice_l118_321) begin
        _zz_when_ArraySlice_l173_321 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_321 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_321 = (_zz_when_ArraySlice_l118_321 <= wReg);
  assign when_ArraySlice_l173_321 = (_zz_when_ArraySlice_l173_321_1 <= _zz_when_ArraySlice_l173_321_3);
  assign when_ArraySlice_l165_322 = (_zz_when_ArraySlice_l165_322 <= selectWriteFifo);
  assign when_ArraySlice_l166_322 = (_zz_when_ArraySlice_l166_322 <= _zz_when_ArraySlice_l166_322_1);
  assign _zz_when_ArraySlice_l112_322 = (wReg % _zz__zz_when_ArraySlice_l112_322);
  assign when_ArraySlice_l112_322 = (_zz_when_ArraySlice_l112_322 != 6'h0);
  assign when_ArraySlice_l113_322 = (7'h40 <= _zz_when_ArraySlice_l113_322);
  always @(*) begin
    if(when_ArraySlice_l112_322) begin
      if(when_ArraySlice_l113_322) begin
        _zz_when_ArraySlice_l173_322 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_322 = (_zz__zz_when_ArraySlice_l173_322 - _zz__zz_when_ArraySlice_l173_322_3);
      end
    end else begin
      if(when_ArraySlice_l118_322) begin
        _zz_when_ArraySlice_l173_322 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_322 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_322 = (_zz_when_ArraySlice_l118_322 <= wReg);
  assign when_ArraySlice_l173_322 = (_zz_when_ArraySlice_l173_322_1 <= _zz_when_ArraySlice_l173_322_3);
  assign when_ArraySlice_l165_323 = (_zz_when_ArraySlice_l165_323 <= selectWriteFifo);
  assign when_ArraySlice_l166_323 = (_zz_when_ArraySlice_l166_323 <= _zz_when_ArraySlice_l166_323_1);
  assign _zz_when_ArraySlice_l112_323 = (wReg % _zz__zz_when_ArraySlice_l112_323);
  assign when_ArraySlice_l112_323 = (_zz_when_ArraySlice_l112_323 != 6'h0);
  assign when_ArraySlice_l113_323 = (7'h40 <= _zz_when_ArraySlice_l113_323);
  always @(*) begin
    if(when_ArraySlice_l112_323) begin
      if(when_ArraySlice_l113_323) begin
        _zz_when_ArraySlice_l173_323 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_323 = (_zz__zz_when_ArraySlice_l173_323 - _zz__zz_when_ArraySlice_l173_323_3);
      end
    end else begin
      if(when_ArraySlice_l118_323) begin
        _zz_when_ArraySlice_l173_323 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_323 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_323 = (_zz_when_ArraySlice_l118_323 <= wReg);
  assign when_ArraySlice_l173_323 = (_zz_when_ArraySlice_l173_323_1 <= _zz_when_ArraySlice_l173_323_3);
  assign when_ArraySlice_l165_324 = (_zz_when_ArraySlice_l165_324 <= selectWriteFifo);
  assign when_ArraySlice_l166_324 = (_zz_when_ArraySlice_l166_324 <= _zz_when_ArraySlice_l166_324_1);
  assign _zz_when_ArraySlice_l112_324 = (wReg % _zz__zz_when_ArraySlice_l112_324);
  assign when_ArraySlice_l112_324 = (_zz_when_ArraySlice_l112_324 != 6'h0);
  assign when_ArraySlice_l113_324 = (7'h40 <= _zz_when_ArraySlice_l113_324);
  always @(*) begin
    if(when_ArraySlice_l112_324) begin
      if(when_ArraySlice_l113_324) begin
        _zz_when_ArraySlice_l173_324 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_324 = (_zz__zz_when_ArraySlice_l173_324 - _zz__zz_when_ArraySlice_l173_324_3);
      end
    end else begin
      if(when_ArraySlice_l118_324) begin
        _zz_when_ArraySlice_l173_324 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_324 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_324 = (_zz_when_ArraySlice_l118_324 <= wReg);
  assign when_ArraySlice_l173_324 = (_zz_when_ArraySlice_l173_324_1 <= _zz_when_ArraySlice_l173_324_3);
  assign when_ArraySlice_l165_325 = (_zz_when_ArraySlice_l165_325 <= selectWriteFifo);
  assign when_ArraySlice_l166_325 = (_zz_when_ArraySlice_l166_325 <= _zz_when_ArraySlice_l166_325_2);
  assign _zz_when_ArraySlice_l112_325 = (wReg % _zz__zz_when_ArraySlice_l112_325);
  assign when_ArraySlice_l112_325 = (_zz_when_ArraySlice_l112_325 != 6'h0);
  assign when_ArraySlice_l113_325 = (7'h40 <= _zz_when_ArraySlice_l113_325);
  always @(*) begin
    if(when_ArraySlice_l112_325) begin
      if(when_ArraySlice_l113_325) begin
        _zz_when_ArraySlice_l173_325 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_325 = (_zz__zz_when_ArraySlice_l173_325 - _zz__zz_when_ArraySlice_l173_325_3);
      end
    end else begin
      if(when_ArraySlice_l118_325) begin
        _zz_when_ArraySlice_l173_325 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_325 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_325 = (_zz_when_ArraySlice_l118_325 <= wReg);
  assign when_ArraySlice_l173_325 = (_zz_when_ArraySlice_l173_325_1 <= _zz_when_ArraySlice_l173_325_3);
  assign when_ArraySlice_l165_326 = (_zz_when_ArraySlice_l165_326 <= selectWriteFifo);
  assign when_ArraySlice_l166_326 = (_zz_when_ArraySlice_l166_326 <= _zz_when_ArraySlice_l166_326_2);
  assign _zz_when_ArraySlice_l112_326 = (wReg % _zz__zz_when_ArraySlice_l112_326);
  assign when_ArraySlice_l112_326 = (_zz_when_ArraySlice_l112_326 != 6'h0);
  assign when_ArraySlice_l113_326 = (7'h40 <= _zz_when_ArraySlice_l113_326);
  always @(*) begin
    if(when_ArraySlice_l112_326) begin
      if(when_ArraySlice_l113_326) begin
        _zz_when_ArraySlice_l173_326 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_326 = (_zz__zz_when_ArraySlice_l173_326 - _zz__zz_when_ArraySlice_l173_326_3);
      end
    end else begin
      if(when_ArraySlice_l118_326) begin
        _zz_when_ArraySlice_l173_326 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_326 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_326 = (_zz_when_ArraySlice_l118_326 <= wReg);
  assign when_ArraySlice_l173_326 = (_zz_when_ArraySlice_l173_326_1 <= _zz_when_ArraySlice_l173_326_3);
  assign when_ArraySlice_l165_327 = (_zz_when_ArraySlice_l165_327 <= selectWriteFifo);
  assign when_ArraySlice_l166_327 = (_zz_when_ArraySlice_l166_327 <= _zz_when_ArraySlice_l166_327_2);
  assign _zz_when_ArraySlice_l112_327 = (wReg % _zz__zz_when_ArraySlice_l112_327);
  assign when_ArraySlice_l112_327 = (_zz_when_ArraySlice_l112_327 != 6'h0);
  assign when_ArraySlice_l113_327 = (7'h40 <= _zz_when_ArraySlice_l113_327);
  always @(*) begin
    if(when_ArraySlice_l112_327) begin
      if(when_ArraySlice_l113_327) begin
        _zz_when_ArraySlice_l173_327 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_327 = (_zz__zz_when_ArraySlice_l173_327 - _zz__zz_when_ArraySlice_l173_327_3);
      end
    end else begin
      if(when_ArraySlice_l118_327) begin
        _zz_when_ArraySlice_l173_327 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_327 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_327 = (_zz_when_ArraySlice_l118_327 <= wReg);
  assign when_ArraySlice_l173_327 = (_zz_when_ArraySlice_l173_327_1 <= _zz_when_ArraySlice_l173_327_3);
  assign when_ArraySlice_l311_4 = (! ((((((_zz_when_ArraySlice_l311_4_1 && _zz_when_ArraySlice_l311_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l311_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l311_4_4 && _zz_when_ArraySlice_l311_4_5) && (debug_4_40 == _zz_when_ArraySlice_l311_4_6)) && (debug_5_40 == 1'b1)) && (debug_6_40 == 1'b1)) && (debug_7_40 == 1'b1))));
  assign outputStreamArrayData_4_fire_12 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l315_4 = ((_zz_when_ArraySlice_l315_4 == 13'h0) && outputStreamArrayData_4_fire_12);
  assign when_ArraySlice_l301_4 = (allowPadding_4 && (wReg <= _zz_when_ArraySlice_l301_4));
  assign outputStreamArrayData_4_fire_13 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l322_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l322_4_1);
  assign when_ArraySlice_l240_5 = (_zz_when_ArraySlice_l240_5 < wReg);
  assign when_ArraySlice_l241_5 = ((! holdReadOp_5) && (_zz_when_ArraySlice_l241_5 != 7'h0));
  assign _zz_outputStreamArrayData_5_valid_1 = (selectReadFifo_5 + _zz__zz_outputStreamArrayData_5_valid_1);
  assign _zz_16 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_5_valid_1);
  assign _zz_io_pop_ready_13 = outputStreamArrayData_5_ready;
  assign when_ArraySlice_l246_5 = (! holdReadOp_5);
  assign outputStreamArrayData_5_fire_7 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l247_5 = ((_zz_when_ArraySlice_l247_5_1 < _zz_when_ArraySlice_l247_5_3) && outputStreamArrayData_5_fire_7);
  assign when_ArraySlice_l248_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l248_5);
  assign when_ArraySlice_l251_5 = (_zz_when_ArraySlice_l251_5 == 13'h0);
  assign outputStreamArrayData_5_fire_8 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l256_5 = ((_zz_when_ArraySlice_l256_5_1 == _zz_when_ArraySlice_l256_5_4) && outputStreamArrayData_5_fire_8);
  assign when_ArraySlice_l257_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l257_5);
  assign _zz_when_ArraySlice_l94_39 = (hReg % _zz__zz_when_ArraySlice_l94_39);
  assign when_ArraySlice_l94_39 = (_zz_when_ArraySlice_l94_39 != 6'h0);
  assign when_ArraySlice_l95_39 = (7'h40 <= _zz_when_ArraySlice_l95_39);
  always @(*) begin
    if(when_ArraySlice_l94_39) begin
      if(when_ArraySlice_l95_39) begin
        _zz_when_ArraySlice_l259_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_5 = (_zz__zz_when_ArraySlice_l259_5 - _zz__zz_when_ArraySlice_l259_5_3);
      end
    end else begin
      if(when_ArraySlice_l99_39) begin
        _zz_when_ArraySlice_l259_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_5 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_39 = (_zz_when_ArraySlice_l99_39 <= hReg);
  assign when_ArraySlice_l259_5 = (_zz_when_ArraySlice_l259_5_1 < _zz_when_ArraySlice_l259_5_4);
  always @(*) begin
    debug_0_41 = 1'b0;
    if(when_ArraySlice_l165_328) begin
      if(when_ArraySlice_l166_328) begin
        debug_0_41 = 1'b1;
      end else begin
        debug_0_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_328) begin
        debug_0_41 = 1'b1;
      end else begin
        debug_0_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_41 = 1'b0;
    if(when_ArraySlice_l165_329) begin
      if(when_ArraySlice_l166_329) begin
        debug_1_41 = 1'b1;
      end else begin
        debug_1_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_329) begin
        debug_1_41 = 1'b1;
      end else begin
        debug_1_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_41 = 1'b0;
    if(when_ArraySlice_l165_330) begin
      if(when_ArraySlice_l166_330) begin
        debug_2_41 = 1'b1;
      end else begin
        debug_2_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_330) begin
        debug_2_41 = 1'b1;
      end else begin
        debug_2_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_41 = 1'b0;
    if(when_ArraySlice_l165_331) begin
      if(when_ArraySlice_l166_331) begin
        debug_3_41 = 1'b1;
      end else begin
        debug_3_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_331) begin
        debug_3_41 = 1'b1;
      end else begin
        debug_3_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_41 = 1'b0;
    if(when_ArraySlice_l165_332) begin
      if(when_ArraySlice_l166_332) begin
        debug_4_41 = 1'b1;
      end else begin
        debug_4_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_332) begin
        debug_4_41 = 1'b1;
      end else begin
        debug_4_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_41 = 1'b0;
    if(when_ArraySlice_l165_333) begin
      if(when_ArraySlice_l166_333) begin
        debug_5_41 = 1'b1;
      end else begin
        debug_5_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_333) begin
        debug_5_41 = 1'b1;
      end else begin
        debug_5_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_41 = 1'b0;
    if(when_ArraySlice_l165_334) begin
      if(when_ArraySlice_l166_334) begin
        debug_6_41 = 1'b1;
      end else begin
        debug_6_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_334) begin
        debug_6_41 = 1'b1;
      end else begin
        debug_6_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_41 = 1'b0;
    if(when_ArraySlice_l165_335) begin
      if(when_ArraySlice_l166_335) begin
        debug_7_41 = 1'b1;
      end else begin
        debug_7_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_335) begin
        debug_7_41 = 1'b1;
      end else begin
        debug_7_41 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_328 = (_zz_when_ArraySlice_l165_328 <= selectWriteFifo);
  assign when_ArraySlice_l166_328 = (_zz_when_ArraySlice_l166_328 <= _zz_when_ArraySlice_l166_328_1);
  assign _zz_when_ArraySlice_l112_328 = (wReg % _zz__zz_when_ArraySlice_l112_328);
  assign when_ArraySlice_l112_328 = (_zz_when_ArraySlice_l112_328 != 6'h0);
  assign when_ArraySlice_l113_328 = (7'h40 <= _zz_when_ArraySlice_l113_328);
  always @(*) begin
    if(when_ArraySlice_l112_328) begin
      if(when_ArraySlice_l113_328) begin
        _zz_when_ArraySlice_l173_328 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_328 = (_zz__zz_when_ArraySlice_l173_328 - _zz__zz_when_ArraySlice_l173_328_3);
      end
    end else begin
      if(when_ArraySlice_l118_328) begin
        _zz_when_ArraySlice_l173_328 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_328 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_328 = (_zz_when_ArraySlice_l118_328 <= wReg);
  assign when_ArraySlice_l173_328 = (_zz_when_ArraySlice_l173_328_1 <= _zz_when_ArraySlice_l173_328_2);
  assign when_ArraySlice_l165_329 = (_zz_when_ArraySlice_l165_329 <= selectWriteFifo);
  assign when_ArraySlice_l166_329 = (_zz_when_ArraySlice_l166_329 <= _zz_when_ArraySlice_l166_329_1);
  assign _zz_when_ArraySlice_l112_329 = (wReg % _zz__zz_when_ArraySlice_l112_329);
  assign when_ArraySlice_l112_329 = (_zz_when_ArraySlice_l112_329 != 6'h0);
  assign when_ArraySlice_l113_329 = (7'h40 <= _zz_when_ArraySlice_l113_329);
  always @(*) begin
    if(when_ArraySlice_l112_329) begin
      if(when_ArraySlice_l113_329) begin
        _zz_when_ArraySlice_l173_329 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_329 = (_zz__zz_when_ArraySlice_l173_329 - _zz__zz_when_ArraySlice_l173_329_3);
      end
    end else begin
      if(when_ArraySlice_l118_329) begin
        _zz_when_ArraySlice_l173_329 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_329 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_329 = (_zz_when_ArraySlice_l118_329 <= wReg);
  assign when_ArraySlice_l173_329 = (_zz_when_ArraySlice_l173_329_1 <= _zz_when_ArraySlice_l173_329_3);
  assign when_ArraySlice_l165_330 = (_zz_when_ArraySlice_l165_330 <= selectWriteFifo);
  assign when_ArraySlice_l166_330 = (_zz_when_ArraySlice_l166_330 <= _zz_when_ArraySlice_l166_330_1);
  assign _zz_when_ArraySlice_l112_330 = (wReg % _zz__zz_when_ArraySlice_l112_330);
  assign when_ArraySlice_l112_330 = (_zz_when_ArraySlice_l112_330 != 6'h0);
  assign when_ArraySlice_l113_330 = (7'h40 <= _zz_when_ArraySlice_l113_330);
  always @(*) begin
    if(when_ArraySlice_l112_330) begin
      if(when_ArraySlice_l113_330) begin
        _zz_when_ArraySlice_l173_330 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_330 = (_zz__zz_when_ArraySlice_l173_330 - _zz__zz_when_ArraySlice_l173_330_3);
      end
    end else begin
      if(when_ArraySlice_l118_330) begin
        _zz_when_ArraySlice_l173_330 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_330 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_330 = (_zz_when_ArraySlice_l118_330 <= wReg);
  assign when_ArraySlice_l173_330 = (_zz_when_ArraySlice_l173_330_1 <= _zz_when_ArraySlice_l173_330_3);
  assign when_ArraySlice_l165_331 = (_zz_when_ArraySlice_l165_331 <= selectWriteFifo);
  assign when_ArraySlice_l166_331 = (_zz_when_ArraySlice_l166_331 <= _zz_when_ArraySlice_l166_331_1);
  assign _zz_when_ArraySlice_l112_331 = (wReg % _zz__zz_when_ArraySlice_l112_331);
  assign when_ArraySlice_l112_331 = (_zz_when_ArraySlice_l112_331 != 6'h0);
  assign when_ArraySlice_l113_331 = (7'h40 <= _zz_when_ArraySlice_l113_331);
  always @(*) begin
    if(when_ArraySlice_l112_331) begin
      if(when_ArraySlice_l113_331) begin
        _zz_when_ArraySlice_l173_331 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_331 = (_zz__zz_when_ArraySlice_l173_331 - _zz__zz_when_ArraySlice_l173_331_3);
      end
    end else begin
      if(when_ArraySlice_l118_331) begin
        _zz_when_ArraySlice_l173_331 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_331 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_331 = (_zz_when_ArraySlice_l118_331 <= wReg);
  assign when_ArraySlice_l173_331 = (_zz_when_ArraySlice_l173_331_1 <= _zz_when_ArraySlice_l173_331_3);
  assign when_ArraySlice_l165_332 = (_zz_when_ArraySlice_l165_332 <= selectWriteFifo);
  assign when_ArraySlice_l166_332 = (_zz_when_ArraySlice_l166_332 <= _zz_when_ArraySlice_l166_332_1);
  assign _zz_when_ArraySlice_l112_332 = (wReg % _zz__zz_when_ArraySlice_l112_332);
  assign when_ArraySlice_l112_332 = (_zz_when_ArraySlice_l112_332 != 6'h0);
  assign when_ArraySlice_l113_332 = (7'h40 <= _zz_when_ArraySlice_l113_332);
  always @(*) begin
    if(when_ArraySlice_l112_332) begin
      if(when_ArraySlice_l113_332) begin
        _zz_when_ArraySlice_l173_332 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_332 = (_zz__zz_when_ArraySlice_l173_332 - _zz__zz_when_ArraySlice_l173_332_3);
      end
    end else begin
      if(when_ArraySlice_l118_332) begin
        _zz_when_ArraySlice_l173_332 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_332 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_332 = (_zz_when_ArraySlice_l118_332 <= wReg);
  assign when_ArraySlice_l173_332 = (_zz_when_ArraySlice_l173_332_1 <= _zz_when_ArraySlice_l173_332_3);
  assign when_ArraySlice_l165_333 = (_zz_when_ArraySlice_l165_333 <= selectWriteFifo);
  assign when_ArraySlice_l166_333 = (_zz_when_ArraySlice_l166_333 <= _zz_when_ArraySlice_l166_333_2);
  assign _zz_when_ArraySlice_l112_333 = (wReg % _zz__zz_when_ArraySlice_l112_333);
  assign when_ArraySlice_l112_333 = (_zz_when_ArraySlice_l112_333 != 6'h0);
  assign when_ArraySlice_l113_333 = (7'h40 <= _zz_when_ArraySlice_l113_333);
  always @(*) begin
    if(when_ArraySlice_l112_333) begin
      if(when_ArraySlice_l113_333) begin
        _zz_when_ArraySlice_l173_333 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_333 = (_zz__zz_when_ArraySlice_l173_333 - _zz__zz_when_ArraySlice_l173_333_3);
      end
    end else begin
      if(when_ArraySlice_l118_333) begin
        _zz_when_ArraySlice_l173_333 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_333 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_333 = (_zz_when_ArraySlice_l118_333 <= wReg);
  assign when_ArraySlice_l173_333 = (_zz_when_ArraySlice_l173_333_1 <= _zz_when_ArraySlice_l173_333_3);
  assign when_ArraySlice_l165_334 = (_zz_when_ArraySlice_l165_334 <= selectWriteFifo);
  assign when_ArraySlice_l166_334 = (_zz_when_ArraySlice_l166_334 <= _zz_when_ArraySlice_l166_334_2);
  assign _zz_when_ArraySlice_l112_334 = (wReg % _zz__zz_when_ArraySlice_l112_334);
  assign when_ArraySlice_l112_334 = (_zz_when_ArraySlice_l112_334 != 6'h0);
  assign when_ArraySlice_l113_334 = (7'h40 <= _zz_when_ArraySlice_l113_334);
  always @(*) begin
    if(when_ArraySlice_l112_334) begin
      if(when_ArraySlice_l113_334) begin
        _zz_when_ArraySlice_l173_334 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_334 = (_zz__zz_when_ArraySlice_l173_334 - _zz__zz_when_ArraySlice_l173_334_3);
      end
    end else begin
      if(when_ArraySlice_l118_334) begin
        _zz_when_ArraySlice_l173_334 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_334 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_334 = (_zz_when_ArraySlice_l118_334 <= wReg);
  assign when_ArraySlice_l173_334 = (_zz_when_ArraySlice_l173_334_1 <= _zz_when_ArraySlice_l173_334_3);
  assign when_ArraySlice_l165_335 = (_zz_when_ArraySlice_l165_335 <= selectWriteFifo);
  assign when_ArraySlice_l166_335 = (_zz_when_ArraySlice_l166_335 <= _zz_when_ArraySlice_l166_335_2);
  assign _zz_when_ArraySlice_l112_335 = (wReg % _zz__zz_when_ArraySlice_l112_335);
  assign when_ArraySlice_l112_335 = (_zz_when_ArraySlice_l112_335 != 6'h0);
  assign when_ArraySlice_l113_335 = (7'h40 <= _zz_when_ArraySlice_l113_335);
  always @(*) begin
    if(when_ArraySlice_l112_335) begin
      if(when_ArraySlice_l113_335) begin
        _zz_when_ArraySlice_l173_335 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_335 = (_zz__zz_when_ArraySlice_l173_335 - _zz__zz_when_ArraySlice_l173_335_3);
      end
    end else begin
      if(when_ArraySlice_l118_335) begin
        _zz_when_ArraySlice_l173_335 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_335 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_335 = (_zz_when_ArraySlice_l118_335 <= wReg);
  assign when_ArraySlice_l173_335 = (_zz_when_ArraySlice_l173_335_1 <= _zz_when_ArraySlice_l173_335_3);
  assign when_ArraySlice_l265_5 = (! ((((((_zz_when_ArraySlice_l265_5_1 && _zz_when_ArraySlice_l265_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l265_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l265_5_4 && _zz_when_ArraySlice_l265_5_5) && (debug_4_41 == _zz_when_ArraySlice_l265_5_6)) && (debug_5_41 == 1'b1)) && (debug_6_41 == 1'b1)) && (debug_7_41 == 1'b1))));
  assign when_ArraySlice_l268_5 = (wReg <= _zz_when_ArraySlice_l268_5_1);
  assign when_ArraySlice_l272_5 = (_zz_when_ArraySlice_l272_5 == 13'h0);
  assign when_ArraySlice_l276_5 = (_zz_when_ArraySlice_l276_5 == 7'h0);
  assign outputStreamArrayData_5_fire_9 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l277_5 = ((handshakeTimes_5_value == _zz_when_ArraySlice_l277_5) && outputStreamArrayData_5_fire_9);
  assign _zz_when_ArraySlice_l94_40 = (hReg % _zz__zz_when_ArraySlice_l94_40);
  assign when_ArraySlice_l94_40 = (_zz_when_ArraySlice_l94_40 != 6'h0);
  assign when_ArraySlice_l95_40 = (7'h40 <= _zz_when_ArraySlice_l95_40);
  always @(*) begin
    if(when_ArraySlice_l94_40) begin
      if(when_ArraySlice_l95_40) begin
        _zz_when_ArraySlice_l279_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_5 = (_zz__zz_when_ArraySlice_l279_5 - _zz__zz_when_ArraySlice_l279_5_3);
      end
    end else begin
      if(when_ArraySlice_l99_40) begin
        _zz_when_ArraySlice_l279_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_5 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_40 = (_zz_when_ArraySlice_l99_40 <= hReg);
  assign when_ArraySlice_l279_5 = (_zz_when_ArraySlice_l279_5_1 < _zz_when_ArraySlice_l279_5_4);
  always @(*) begin
    debug_0_42 = 1'b0;
    if(when_ArraySlice_l165_336) begin
      if(when_ArraySlice_l166_336) begin
        debug_0_42 = 1'b1;
      end else begin
        debug_0_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_336) begin
        debug_0_42 = 1'b1;
      end else begin
        debug_0_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_42 = 1'b0;
    if(when_ArraySlice_l165_337) begin
      if(when_ArraySlice_l166_337) begin
        debug_1_42 = 1'b1;
      end else begin
        debug_1_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_337) begin
        debug_1_42 = 1'b1;
      end else begin
        debug_1_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_42 = 1'b0;
    if(when_ArraySlice_l165_338) begin
      if(when_ArraySlice_l166_338) begin
        debug_2_42 = 1'b1;
      end else begin
        debug_2_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_338) begin
        debug_2_42 = 1'b1;
      end else begin
        debug_2_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_42 = 1'b0;
    if(when_ArraySlice_l165_339) begin
      if(when_ArraySlice_l166_339) begin
        debug_3_42 = 1'b1;
      end else begin
        debug_3_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_339) begin
        debug_3_42 = 1'b1;
      end else begin
        debug_3_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_42 = 1'b0;
    if(when_ArraySlice_l165_340) begin
      if(when_ArraySlice_l166_340) begin
        debug_4_42 = 1'b1;
      end else begin
        debug_4_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_340) begin
        debug_4_42 = 1'b1;
      end else begin
        debug_4_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_42 = 1'b0;
    if(when_ArraySlice_l165_341) begin
      if(when_ArraySlice_l166_341) begin
        debug_5_42 = 1'b1;
      end else begin
        debug_5_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_341) begin
        debug_5_42 = 1'b1;
      end else begin
        debug_5_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_42 = 1'b0;
    if(when_ArraySlice_l165_342) begin
      if(when_ArraySlice_l166_342) begin
        debug_6_42 = 1'b1;
      end else begin
        debug_6_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_342) begin
        debug_6_42 = 1'b1;
      end else begin
        debug_6_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_42 = 1'b0;
    if(when_ArraySlice_l165_343) begin
      if(when_ArraySlice_l166_343) begin
        debug_7_42 = 1'b1;
      end else begin
        debug_7_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_343) begin
        debug_7_42 = 1'b1;
      end else begin
        debug_7_42 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_336 = (_zz_when_ArraySlice_l165_336 <= selectWriteFifo);
  assign when_ArraySlice_l166_336 = (_zz_when_ArraySlice_l166_336 <= _zz_when_ArraySlice_l166_336_1);
  assign _zz_when_ArraySlice_l112_336 = (wReg % _zz__zz_when_ArraySlice_l112_336);
  assign when_ArraySlice_l112_336 = (_zz_when_ArraySlice_l112_336 != 6'h0);
  assign when_ArraySlice_l113_336 = (7'h40 <= _zz_when_ArraySlice_l113_336);
  always @(*) begin
    if(when_ArraySlice_l112_336) begin
      if(when_ArraySlice_l113_336) begin
        _zz_when_ArraySlice_l173_336 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_336 = (_zz__zz_when_ArraySlice_l173_336 - _zz__zz_when_ArraySlice_l173_336_3);
      end
    end else begin
      if(when_ArraySlice_l118_336) begin
        _zz_when_ArraySlice_l173_336 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_336 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_336 = (_zz_when_ArraySlice_l118_336 <= wReg);
  assign when_ArraySlice_l173_336 = (_zz_when_ArraySlice_l173_336_1 <= _zz_when_ArraySlice_l173_336_2);
  assign when_ArraySlice_l165_337 = (_zz_when_ArraySlice_l165_337 <= selectWriteFifo);
  assign when_ArraySlice_l166_337 = (_zz_when_ArraySlice_l166_337 <= _zz_when_ArraySlice_l166_337_1);
  assign _zz_when_ArraySlice_l112_337 = (wReg % _zz__zz_when_ArraySlice_l112_337);
  assign when_ArraySlice_l112_337 = (_zz_when_ArraySlice_l112_337 != 6'h0);
  assign when_ArraySlice_l113_337 = (7'h40 <= _zz_when_ArraySlice_l113_337);
  always @(*) begin
    if(when_ArraySlice_l112_337) begin
      if(when_ArraySlice_l113_337) begin
        _zz_when_ArraySlice_l173_337 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_337 = (_zz__zz_when_ArraySlice_l173_337 - _zz__zz_when_ArraySlice_l173_337_3);
      end
    end else begin
      if(when_ArraySlice_l118_337) begin
        _zz_when_ArraySlice_l173_337 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_337 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_337 = (_zz_when_ArraySlice_l118_337 <= wReg);
  assign when_ArraySlice_l173_337 = (_zz_when_ArraySlice_l173_337_1 <= _zz_when_ArraySlice_l173_337_3);
  assign when_ArraySlice_l165_338 = (_zz_when_ArraySlice_l165_338 <= selectWriteFifo);
  assign when_ArraySlice_l166_338 = (_zz_when_ArraySlice_l166_338 <= _zz_when_ArraySlice_l166_338_1);
  assign _zz_when_ArraySlice_l112_338 = (wReg % _zz__zz_when_ArraySlice_l112_338);
  assign when_ArraySlice_l112_338 = (_zz_when_ArraySlice_l112_338 != 6'h0);
  assign when_ArraySlice_l113_338 = (7'h40 <= _zz_when_ArraySlice_l113_338);
  always @(*) begin
    if(when_ArraySlice_l112_338) begin
      if(when_ArraySlice_l113_338) begin
        _zz_when_ArraySlice_l173_338 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_338 = (_zz__zz_when_ArraySlice_l173_338 - _zz__zz_when_ArraySlice_l173_338_3);
      end
    end else begin
      if(when_ArraySlice_l118_338) begin
        _zz_when_ArraySlice_l173_338 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_338 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_338 = (_zz_when_ArraySlice_l118_338 <= wReg);
  assign when_ArraySlice_l173_338 = (_zz_when_ArraySlice_l173_338_1 <= _zz_when_ArraySlice_l173_338_3);
  assign when_ArraySlice_l165_339 = (_zz_when_ArraySlice_l165_339 <= selectWriteFifo);
  assign when_ArraySlice_l166_339 = (_zz_when_ArraySlice_l166_339 <= _zz_when_ArraySlice_l166_339_1);
  assign _zz_when_ArraySlice_l112_339 = (wReg % _zz__zz_when_ArraySlice_l112_339);
  assign when_ArraySlice_l112_339 = (_zz_when_ArraySlice_l112_339 != 6'h0);
  assign when_ArraySlice_l113_339 = (7'h40 <= _zz_when_ArraySlice_l113_339);
  always @(*) begin
    if(when_ArraySlice_l112_339) begin
      if(when_ArraySlice_l113_339) begin
        _zz_when_ArraySlice_l173_339 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_339 = (_zz__zz_when_ArraySlice_l173_339 - _zz__zz_when_ArraySlice_l173_339_3);
      end
    end else begin
      if(when_ArraySlice_l118_339) begin
        _zz_when_ArraySlice_l173_339 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_339 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_339 = (_zz_when_ArraySlice_l118_339 <= wReg);
  assign when_ArraySlice_l173_339 = (_zz_when_ArraySlice_l173_339_1 <= _zz_when_ArraySlice_l173_339_3);
  assign when_ArraySlice_l165_340 = (_zz_when_ArraySlice_l165_340 <= selectWriteFifo);
  assign when_ArraySlice_l166_340 = (_zz_when_ArraySlice_l166_340 <= _zz_when_ArraySlice_l166_340_1);
  assign _zz_when_ArraySlice_l112_340 = (wReg % _zz__zz_when_ArraySlice_l112_340);
  assign when_ArraySlice_l112_340 = (_zz_when_ArraySlice_l112_340 != 6'h0);
  assign when_ArraySlice_l113_340 = (7'h40 <= _zz_when_ArraySlice_l113_340);
  always @(*) begin
    if(when_ArraySlice_l112_340) begin
      if(when_ArraySlice_l113_340) begin
        _zz_when_ArraySlice_l173_340 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_340 = (_zz__zz_when_ArraySlice_l173_340 - _zz__zz_when_ArraySlice_l173_340_3);
      end
    end else begin
      if(when_ArraySlice_l118_340) begin
        _zz_when_ArraySlice_l173_340 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_340 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_340 = (_zz_when_ArraySlice_l118_340 <= wReg);
  assign when_ArraySlice_l173_340 = (_zz_when_ArraySlice_l173_340_1 <= _zz_when_ArraySlice_l173_340_3);
  assign when_ArraySlice_l165_341 = (_zz_when_ArraySlice_l165_341 <= selectWriteFifo);
  assign when_ArraySlice_l166_341 = (_zz_when_ArraySlice_l166_341 <= _zz_when_ArraySlice_l166_341_2);
  assign _zz_when_ArraySlice_l112_341 = (wReg % _zz__zz_when_ArraySlice_l112_341);
  assign when_ArraySlice_l112_341 = (_zz_when_ArraySlice_l112_341 != 6'h0);
  assign when_ArraySlice_l113_341 = (7'h40 <= _zz_when_ArraySlice_l113_341);
  always @(*) begin
    if(when_ArraySlice_l112_341) begin
      if(when_ArraySlice_l113_341) begin
        _zz_when_ArraySlice_l173_341 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_341 = (_zz__zz_when_ArraySlice_l173_341 - _zz__zz_when_ArraySlice_l173_341_3);
      end
    end else begin
      if(when_ArraySlice_l118_341) begin
        _zz_when_ArraySlice_l173_341 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_341 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_341 = (_zz_when_ArraySlice_l118_341 <= wReg);
  assign when_ArraySlice_l173_341 = (_zz_when_ArraySlice_l173_341_1 <= _zz_when_ArraySlice_l173_341_3);
  assign when_ArraySlice_l165_342 = (_zz_when_ArraySlice_l165_342 <= selectWriteFifo);
  assign when_ArraySlice_l166_342 = (_zz_when_ArraySlice_l166_342 <= _zz_when_ArraySlice_l166_342_2);
  assign _zz_when_ArraySlice_l112_342 = (wReg % _zz__zz_when_ArraySlice_l112_342);
  assign when_ArraySlice_l112_342 = (_zz_when_ArraySlice_l112_342 != 6'h0);
  assign when_ArraySlice_l113_342 = (7'h40 <= _zz_when_ArraySlice_l113_342);
  always @(*) begin
    if(when_ArraySlice_l112_342) begin
      if(when_ArraySlice_l113_342) begin
        _zz_when_ArraySlice_l173_342 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_342 = (_zz__zz_when_ArraySlice_l173_342 - _zz__zz_when_ArraySlice_l173_342_3);
      end
    end else begin
      if(when_ArraySlice_l118_342) begin
        _zz_when_ArraySlice_l173_342 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_342 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_342 = (_zz_when_ArraySlice_l118_342 <= wReg);
  assign when_ArraySlice_l173_342 = (_zz_when_ArraySlice_l173_342_1 <= _zz_when_ArraySlice_l173_342_3);
  assign when_ArraySlice_l165_343 = (_zz_when_ArraySlice_l165_343 <= selectWriteFifo);
  assign when_ArraySlice_l166_343 = (_zz_when_ArraySlice_l166_343 <= _zz_when_ArraySlice_l166_343_2);
  assign _zz_when_ArraySlice_l112_343 = (wReg % _zz__zz_when_ArraySlice_l112_343);
  assign when_ArraySlice_l112_343 = (_zz_when_ArraySlice_l112_343 != 6'h0);
  assign when_ArraySlice_l113_343 = (7'h40 <= _zz_when_ArraySlice_l113_343);
  always @(*) begin
    if(when_ArraySlice_l112_343) begin
      if(when_ArraySlice_l113_343) begin
        _zz_when_ArraySlice_l173_343 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_343 = (_zz__zz_when_ArraySlice_l173_343 - _zz__zz_when_ArraySlice_l173_343_3);
      end
    end else begin
      if(when_ArraySlice_l118_343) begin
        _zz_when_ArraySlice_l173_343 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_343 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_343 = (_zz_when_ArraySlice_l118_343 <= wReg);
  assign when_ArraySlice_l173_343 = (_zz_when_ArraySlice_l173_343_1 <= _zz_when_ArraySlice_l173_343_3);
  assign when_ArraySlice_l285_5 = (! ((((((_zz_when_ArraySlice_l285_5_1 && _zz_when_ArraySlice_l285_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l285_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l285_5_4 && _zz_when_ArraySlice_l285_5_5) && (debug_4_42 == _zz_when_ArraySlice_l285_5_6)) && (debug_5_42 == 1'b1)) && (debug_6_42 == 1'b1)) && (debug_7_42 == 1'b1))));
  assign when_ArraySlice_l288_5 = (wReg <= _zz_when_ArraySlice_l288_5_1);
  assign outputStreamArrayData_5_fire_10 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l292_5 = ((_zz_when_ArraySlice_l292_5 == 13'h0) && outputStreamArrayData_5_fire_10);
  assign outputStreamArrayData_5_fire_11 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l303_5 = ((handshakeTimes_5_value == _zz_when_ArraySlice_l303_5) && outputStreamArrayData_5_fire_11);
  assign _zz_when_ArraySlice_l94_41 = (hReg % _zz__zz_when_ArraySlice_l94_41);
  assign when_ArraySlice_l94_41 = (_zz_when_ArraySlice_l94_41 != 6'h0);
  assign when_ArraySlice_l95_41 = (7'h40 <= _zz_when_ArraySlice_l95_41);
  always @(*) begin
    if(when_ArraySlice_l94_41) begin
      if(when_ArraySlice_l95_41) begin
        _zz_when_ArraySlice_l304_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_5 = (_zz__zz_when_ArraySlice_l304_5 - _zz__zz_when_ArraySlice_l304_5_3);
      end
    end else begin
      if(when_ArraySlice_l99_41) begin
        _zz_when_ArraySlice_l304_5 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_5 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_41 = (_zz_when_ArraySlice_l99_41 <= hReg);
  assign when_ArraySlice_l304_5 = (_zz_when_ArraySlice_l304_5_1 < _zz_when_ArraySlice_l304_5_4);
  always @(*) begin
    debug_0_43 = 1'b0;
    if(when_ArraySlice_l165_344) begin
      if(when_ArraySlice_l166_344) begin
        debug_0_43 = 1'b1;
      end else begin
        debug_0_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_344) begin
        debug_0_43 = 1'b1;
      end else begin
        debug_0_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_43 = 1'b0;
    if(when_ArraySlice_l165_345) begin
      if(when_ArraySlice_l166_345) begin
        debug_1_43 = 1'b1;
      end else begin
        debug_1_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_345) begin
        debug_1_43 = 1'b1;
      end else begin
        debug_1_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_43 = 1'b0;
    if(when_ArraySlice_l165_346) begin
      if(when_ArraySlice_l166_346) begin
        debug_2_43 = 1'b1;
      end else begin
        debug_2_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_346) begin
        debug_2_43 = 1'b1;
      end else begin
        debug_2_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_43 = 1'b0;
    if(when_ArraySlice_l165_347) begin
      if(when_ArraySlice_l166_347) begin
        debug_3_43 = 1'b1;
      end else begin
        debug_3_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_347) begin
        debug_3_43 = 1'b1;
      end else begin
        debug_3_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_43 = 1'b0;
    if(when_ArraySlice_l165_348) begin
      if(when_ArraySlice_l166_348) begin
        debug_4_43 = 1'b1;
      end else begin
        debug_4_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_348) begin
        debug_4_43 = 1'b1;
      end else begin
        debug_4_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_43 = 1'b0;
    if(when_ArraySlice_l165_349) begin
      if(when_ArraySlice_l166_349) begin
        debug_5_43 = 1'b1;
      end else begin
        debug_5_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_349) begin
        debug_5_43 = 1'b1;
      end else begin
        debug_5_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_43 = 1'b0;
    if(when_ArraySlice_l165_350) begin
      if(when_ArraySlice_l166_350) begin
        debug_6_43 = 1'b1;
      end else begin
        debug_6_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_350) begin
        debug_6_43 = 1'b1;
      end else begin
        debug_6_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_43 = 1'b0;
    if(when_ArraySlice_l165_351) begin
      if(when_ArraySlice_l166_351) begin
        debug_7_43 = 1'b1;
      end else begin
        debug_7_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_351) begin
        debug_7_43 = 1'b1;
      end else begin
        debug_7_43 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_344 = (_zz_when_ArraySlice_l165_344 <= selectWriteFifo);
  assign when_ArraySlice_l166_344 = (_zz_when_ArraySlice_l166_344 <= _zz_when_ArraySlice_l166_344_1);
  assign _zz_when_ArraySlice_l112_344 = (wReg % _zz__zz_when_ArraySlice_l112_344);
  assign when_ArraySlice_l112_344 = (_zz_when_ArraySlice_l112_344 != 6'h0);
  assign when_ArraySlice_l113_344 = (7'h40 <= _zz_when_ArraySlice_l113_344);
  always @(*) begin
    if(when_ArraySlice_l112_344) begin
      if(when_ArraySlice_l113_344) begin
        _zz_when_ArraySlice_l173_344 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_344 = (_zz__zz_when_ArraySlice_l173_344 - _zz__zz_when_ArraySlice_l173_344_3);
      end
    end else begin
      if(when_ArraySlice_l118_344) begin
        _zz_when_ArraySlice_l173_344 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_344 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_344 = (_zz_when_ArraySlice_l118_344 <= wReg);
  assign when_ArraySlice_l173_344 = (_zz_when_ArraySlice_l173_344_1 <= _zz_when_ArraySlice_l173_344_2);
  assign when_ArraySlice_l165_345 = (_zz_when_ArraySlice_l165_345 <= selectWriteFifo);
  assign when_ArraySlice_l166_345 = (_zz_when_ArraySlice_l166_345 <= _zz_when_ArraySlice_l166_345_1);
  assign _zz_when_ArraySlice_l112_345 = (wReg % _zz__zz_when_ArraySlice_l112_345);
  assign when_ArraySlice_l112_345 = (_zz_when_ArraySlice_l112_345 != 6'h0);
  assign when_ArraySlice_l113_345 = (7'h40 <= _zz_when_ArraySlice_l113_345);
  always @(*) begin
    if(when_ArraySlice_l112_345) begin
      if(when_ArraySlice_l113_345) begin
        _zz_when_ArraySlice_l173_345 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_345 = (_zz__zz_when_ArraySlice_l173_345 - _zz__zz_when_ArraySlice_l173_345_3);
      end
    end else begin
      if(when_ArraySlice_l118_345) begin
        _zz_when_ArraySlice_l173_345 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_345 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_345 = (_zz_when_ArraySlice_l118_345 <= wReg);
  assign when_ArraySlice_l173_345 = (_zz_when_ArraySlice_l173_345_1 <= _zz_when_ArraySlice_l173_345_3);
  assign when_ArraySlice_l165_346 = (_zz_when_ArraySlice_l165_346 <= selectWriteFifo);
  assign when_ArraySlice_l166_346 = (_zz_when_ArraySlice_l166_346 <= _zz_when_ArraySlice_l166_346_1);
  assign _zz_when_ArraySlice_l112_346 = (wReg % _zz__zz_when_ArraySlice_l112_346);
  assign when_ArraySlice_l112_346 = (_zz_when_ArraySlice_l112_346 != 6'h0);
  assign when_ArraySlice_l113_346 = (7'h40 <= _zz_when_ArraySlice_l113_346);
  always @(*) begin
    if(when_ArraySlice_l112_346) begin
      if(when_ArraySlice_l113_346) begin
        _zz_when_ArraySlice_l173_346 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_346 = (_zz__zz_when_ArraySlice_l173_346 - _zz__zz_when_ArraySlice_l173_346_3);
      end
    end else begin
      if(when_ArraySlice_l118_346) begin
        _zz_when_ArraySlice_l173_346 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_346 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_346 = (_zz_when_ArraySlice_l118_346 <= wReg);
  assign when_ArraySlice_l173_346 = (_zz_when_ArraySlice_l173_346_1 <= _zz_when_ArraySlice_l173_346_3);
  assign when_ArraySlice_l165_347 = (_zz_when_ArraySlice_l165_347 <= selectWriteFifo);
  assign when_ArraySlice_l166_347 = (_zz_when_ArraySlice_l166_347 <= _zz_when_ArraySlice_l166_347_1);
  assign _zz_when_ArraySlice_l112_347 = (wReg % _zz__zz_when_ArraySlice_l112_347);
  assign when_ArraySlice_l112_347 = (_zz_when_ArraySlice_l112_347 != 6'h0);
  assign when_ArraySlice_l113_347 = (7'h40 <= _zz_when_ArraySlice_l113_347);
  always @(*) begin
    if(when_ArraySlice_l112_347) begin
      if(when_ArraySlice_l113_347) begin
        _zz_when_ArraySlice_l173_347 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_347 = (_zz__zz_when_ArraySlice_l173_347 - _zz__zz_when_ArraySlice_l173_347_3);
      end
    end else begin
      if(when_ArraySlice_l118_347) begin
        _zz_when_ArraySlice_l173_347 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_347 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_347 = (_zz_when_ArraySlice_l118_347 <= wReg);
  assign when_ArraySlice_l173_347 = (_zz_when_ArraySlice_l173_347_1 <= _zz_when_ArraySlice_l173_347_3);
  assign when_ArraySlice_l165_348 = (_zz_when_ArraySlice_l165_348 <= selectWriteFifo);
  assign when_ArraySlice_l166_348 = (_zz_when_ArraySlice_l166_348 <= _zz_when_ArraySlice_l166_348_1);
  assign _zz_when_ArraySlice_l112_348 = (wReg % _zz__zz_when_ArraySlice_l112_348);
  assign when_ArraySlice_l112_348 = (_zz_when_ArraySlice_l112_348 != 6'h0);
  assign when_ArraySlice_l113_348 = (7'h40 <= _zz_when_ArraySlice_l113_348);
  always @(*) begin
    if(when_ArraySlice_l112_348) begin
      if(when_ArraySlice_l113_348) begin
        _zz_when_ArraySlice_l173_348 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_348 = (_zz__zz_when_ArraySlice_l173_348 - _zz__zz_when_ArraySlice_l173_348_3);
      end
    end else begin
      if(when_ArraySlice_l118_348) begin
        _zz_when_ArraySlice_l173_348 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_348 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_348 = (_zz_when_ArraySlice_l118_348 <= wReg);
  assign when_ArraySlice_l173_348 = (_zz_when_ArraySlice_l173_348_1 <= _zz_when_ArraySlice_l173_348_3);
  assign when_ArraySlice_l165_349 = (_zz_when_ArraySlice_l165_349 <= selectWriteFifo);
  assign when_ArraySlice_l166_349 = (_zz_when_ArraySlice_l166_349 <= _zz_when_ArraySlice_l166_349_2);
  assign _zz_when_ArraySlice_l112_349 = (wReg % _zz__zz_when_ArraySlice_l112_349);
  assign when_ArraySlice_l112_349 = (_zz_when_ArraySlice_l112_349 != 6'h0);
  assign when_ArraySlice_l113_349 = (7'h40 <= _zz_when_ArraySlice_l113_349);
  always @(*) begin
    if(when_ArraySlice_l112_349) begin
      if(when_ArraySlice_l113_349) begin
        _zz_when_ArraySlice_l173_349 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_349 = (_zz__zz_when_ArraySlice_l173_349 - _zz__zz_when_ArraySlice_l173_349_3);
      end
    end else begin
      if(when_ArraySlice_l118_349) begin
        _zz_when_ArraySlice_l173_349 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_349 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_349 = (_zz_when_ArraySlice_l118_349 <= wReg);
  assign when_ArraySlice_l173_349 = (_zz_when_ArraySlice_l173_349_1 <= _zz_when_ArraySlice_l173_349_3);
  assign when_ArraySlice_l165_350 = (_zz_when_ArraySlice_l165_350 <= selectWriteFifo);
  assign when_ArraySlice_l166_350 = (_zz_when_ArraySlice_l166_350 <= _zz_when_ArraySlice_l166_350_2);
  assign _zz_when_ArraySlice_l112_350 = (wReg % _zz__zz_when_ArraySlice_l112_350);
  assign when_ArraySlice_l112_350 = (_zz_when_ArraySlice_l112_350 != 6'h0);
  assign when_ArraySlice_l113_350 = (7'h40 <= _zz_when_ArraySlice_l113_350);
  always @(*) begin
    if(when_ArraySlice_l112_350) begin
      if(when_ArraySlice_l113_350) begin
        _zz_when_ArraySlice_l173_350 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_350 = (_zz__zz_when_ArraySlice_l173_350 - _zz__zz_when_ArraySlice_l173_350_3);
      end
    end else begin
      if(when_ArraySlice_l118_350) begin
        _zz_when_ArraySlice_l173_350 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_350 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_350 = (_zz_when_ArraySlice_l118_350 <= wReg);
  assign when_ArraySlice_l173_350 = (_zz_when_ArraySlice_l173_350_1 <= _zz_when_ArraySlice_l173_350_3);
  assign when_ArraySlice_l165_351 = (_zz_when_ArraySlice_l165_351 <= selectWriteFifo);
  assign when_ArraySlice_l166_351 = (_zz_when_ArraySlice_l166_351 <= _zz_when_ArraySlice_l166_351_2);
  assign _zz_when_ArraySlice_l112_351 = (wReg % _zz__zz_when_ArraySlice_l112_351);
  assign when_ArraySlice_l112_351 = (_zz_when_ArraySlice_l112_351 != 6'h0);
  assign when_ArraySlice_l113_351 = (7'h40 <= _zz_when_ArraySlice_l113_351);
  always @(*) begin
    if(when_ArraySlice_l112_351) begin
      if(when_ArraySlice_l113_351) begin
        _zz_when_ArraySlice_l173_351 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_351 = (_zz__zz_when_ArraySlice_l173_351 - _zz__zz_when_ArraySlice_l173_351_3);
      end
    end else begin
      if(when_ArraySlice_l118_351) begin
        _zz_when_ArraySlice_l173_351 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_351 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_351 = (_zz_when_ArraySlice_l118_351 <= wReg);
  assign when_ArraySlice_l173_351 = (_zz_when_ArraySlice_l173_351_1 <= _zz_when_ArraySlice_l173_351_3);
  assign when_ArraySlice_l311_5 = (! ((((((_zz_when_ArraySlice_l311_5_1 && _zz_when_ArraySlice_l311_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l311_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l311_5_4 && _zz_when_ArraySlice_l311_5_5) && (debug_4_43 == _zz_when_ArraySlice_l311_5_6)) && (debug_5_43 == 1'b1)) && (debug_6_43 == 1'b1)) && (debug_7_43 == 1'b1))));
  assign outputStreamArrayData_5_fire_12 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l315_5 = ((_zz_when_ArraySlice_l315_5 == 13'h0) && outputStreamArrayData_5_fire_12);
  assign when_ArraySlice_l301_5 = (allowPadding_5 && (wReg <= _zz_when_ArraySlice_l301_5));
  assign outputStreamArrayData_5_fire_13 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l322_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l322_5);
  assign when_ArraySlice_l240_6 = (_zz_when_ArraySlice_l240_6 < wReg);
  assign when_ArraySlice_l241_6 = ((! holdReadOp_6) && (_zz_when_ArraySlice_l241_6 != 7'h0));
  assign _zz_outputStreamArrayData_6_valid_1 = (selectReadFifo_6 + _zz__zz_outputStreamArrayData_6_valid_1);
  assign _zz_17 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_6_valid_1);
  assign _zz_io_pop_ready_14 = outputStreamArrayData_6_ready;
  assign when_ArraySlice_l246_6 = (! holdReadOp_6);
  assign outputStreamArrayData_6_fire_7 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l247_6 = ((_zz_when_ArraySlice_l247_6 < _zz_when_ArraySlice_l247_6_2) && outputStreamArrayData_6_fire_7);
  assign when_ArraySlice_l248_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l248_6);
  assign when_ArraySlice_l251_6 = (_zz_when_ArraySlice_l251_6 == 13'h0);
  assign outputStreamArrayData_6_fire_8 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l256_6 = ((_zz_when_ArraySlice_l256_6 == _zz_when_ArraySlice_l256_6_3) && outputStreamArrayData_6_fire_8);
  assign when_ArraySlice_l257_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l257_6);
  assign _zz_when_ArraySlice_l94_42 = (hReg % _zz__zz_when_ArraySlice_l94_42);
  assign when_ArraySlice_l94_42 = (_zz_when_ArraySlice_l94_42 != 6'h0);
  assign when_ArraySlice_l95_42 = (7'h40 <= _zz_when_ArraySlice_l95_42);
  always @(*) begin
    if(when_ArraySlice_l94_42) begin
      if(when_ArraySlice_l95_42) begin
        _zz_when_ArraySlice_l259_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_6 = (_zz__zz_when_ArraySlice_l259_6 - _zz__zz_when_ArraySlice_l259_6_3);
      end
    end else begin
      if(when_ArraySlice_l99_42) begin
        _zz_when_ArraySlice_l259_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_6 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_42 = (_zz_when_ArraySlice_l99_42 <= hReg);
  assign when_ArraySlice_l259_6 = (_zz_when_ArraySlice_l259_6_1 < _zz_when_ArraySlice_l259_6_4);
  always @(*) begin
    debug_0_44 = 1'b0;
    if(when_ArraySlice_l165_352) begin
      if(when_ArraySlice_l166_352) begin
        debug_0_44 = 1'b1;
      end else begin
        debug_0_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_352) begin
        debug_0_44 = 1'b1;
      end else begin
        debug_0_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_44 = 1'b0;
    if(when_ArraySlice_l165_353) begin
      if(when_ArraySlice_l166_353) begin
        debug_1_44 = 1'b1;
      end else begin
        debug_1_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_353) begin
        debug_1_44 = 1'b1;
      end else begin
        debug_1_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_44 = 1'b0;
    if(when_ArraySlice_l165_354) begin
      if(when_ArraySlice_l166_354) begin
        debug_2_44 = 1'b1;
      end else begin
        debug_2_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_354) begin
        debug_2_44 = 1'b1;
      end else begin
        debug_2_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_44 = 1'b0;
    if(when_ArraySlice_l165_355) begin
      if(when_ArraySlice_l166_355) begin
        debug_3_44 = 1'b1;
      end else begin
        debug_3_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_355) begin
        debug_3_44 = 1'b1;
      end else begin
        debug_3_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_44 = 1'b0;
    if(when_ArraySlice_l165_356) begin
      if(when_ArraySlice_l166_356) begin
        debug_4_44 = 1'b1;
      end else begin
        debug_4_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_356) begin
        debug_4_44 = 1'b1;
      end else begin
        debug_4_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_44 = 1'b0;
    if(when_ArraySlice_l165_357) begin
      if(when_ArraySlice_l166_357) begin
        debug_5_44 = 1'b1;
      end else begin
        debug_5_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_357) begin
        debug_5_44 = 1'b1;
      end else begin
        debug_5_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_44 = 1'b0;
    if(when_ArraySlice_l165_358) begin
      if(when_ArraySlice_l166_358) begin
        debug_6_44 = 1'b1;
      end else begin
        debug_6_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_358) begin
        debug_6_44 = 1'b1;
      end else begin
        debug_6_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_44 = 1'b0;
    if(when_ArraySlice_l165_359) begin
      if(when_ArraySlice_l166_359) begin
        debug_7_44 = 1'b1;
      end else begin
        debug_7_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_359) begin
        debug_7_44 = 1'b1;
      end else begin
        debug_7_44 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_352 = (_zz_when_ArraySlice_l165_352 <= selectWriteFifo);
  assign when_ArraySlice_l166_352 = (_zz_when_ArraySlice_l166_352 <= _zz_when_ArraySlice_l166_352_1);
  assign _zz_when_ArraySlice_l112_352 = (wReg % _zz__zz_when_ArraySlice_l112_352);
  assign when_ArraySlice_l112_352 = (_zz_when_ArraySlice_l112_352 != 6'h0);
  assign when_ArraySlice_l113_352 = (7'h40 <= _zz_when_ArraySlice_l113_352);
  always @(*) begin
    if(when_ArraySlice_l112_352) begin
      if(when_ArraySlice_l113_352) begin
        _zz_when_ArraySlice_l173_352 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_352 = (_zz__zz_when_ArraySlice_l173_352 - _zz__zz_when_ArraySlice_l173_352_3);
      end
    end else begin
      if(when_ArraySlice_l118_352) begin
        _zz_when_ArraySlice_l173_352 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_352 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_352 = (_zz_when_ArraySlice_l118_352 <= wReg);
  assign when_ArraySlice_l173_352 = (_zz_when_ArraySlice_l173_352_1 <= _zz_when_ArraySlice_l173_352_2);
  assign when_ArraySlice_l165_353 = (_zz_when_ArraySlice_l165_353 <= selectWriteFifo);
  assign when_ArraySlice_l166_353 = (_zz_when_ArraySlice_l166_353 <= _zz_when_ArraySlice_l166_353_1);
  assign _zz_when_ArraySlice_l112_353 = (wReg % _zz__zz_when_ArraySlice_l112_353);
  assign when_ArraySlice_l112_353 = (_zz_when_ArraySlice_l112_353 != 6'h0);
  assign when_ArraySlice_l113_353 = (7'h40 <= _zz_when_ArraySlice_l113_353);
  always @(*) begin
    if(when_ArraySlice_l112_353) begin
      if(when_ArraySlice_l113_353) begin
        _zz_when_ArraySlice_l173_353 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_353 = (_zz__zz_when_ArraySlice_l173_353 - _zz__zz_when_ArraySlice_l173_353_3);
      end
    end else begin
      if(when_ArraySlice_l118_353) begin
        _zz_when_ArraySlice_l173_353 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_353 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_353 = (_zz_when_ArraySlice_l118_353 <= wReg);
  assign when_ArraySlice_l173_353 = (_zz_when_ArraySlice_l173_353_1 <= _zz_when_ArraySlice_l173_353_3);
  assign when_ArraySlice_l165_354 = (_zz_when_ArraySlice_l165_354 <= selectWriteFifo);
  assign when_ArraySlice_l166_354 = (_zz_when_ArraySlice_l166_354 <= _zz_when_ArraySlice_l166_354_1);
  assign _zz_when_ArraySlice_l112_354 = (wReg % _zz__zz_when_ArraySlice_l112_354);
  assign when_ArraySlice_l112_354 = (_zz_when_ArraySlice_l112_354 != 6'h0);
  assign when_ArraySlice_l113_354 = (7'h40 <= _zz_when_ArraySlice_l113_354);
  always @(*) begin
    if(when_ArraySlice_l112_354) begin
      if(when_ArraySlice_l113_354) begin
        _zz_when_ArraySlice_l173_354 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_354 = (_zz__zz_when_ArraySlice_l173_354 - _zz__zz_when_ArraySlice_l173_354_3);
      end
    end else begin
      if(when_ArraySlice_l118_354) begin
        _zz_when_ArraySlice_l173_354 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_354 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_354 = (_zz_when_ArraySlice_l118_354 <= wReg);
  assign when_ArraySlice_l173_354 = (_zz_when_ArraySlice_l173_354_1 <= _zz_when_ArraySlice_l173_354_3);
  assign when_ArraySlice_l165_355 = (_zz_when_ArraySlice_l165_355 <= selectWriteFifo);
  assign when_ArraySlice_l166_355 = (_zz_when_ArraySlice_l166_355 <= _zz_when_ArraySlice_l166_355_1);
  assign _zz_when_ArraySlice_l112_355 = (wReg % _zz__zz_when_ArraySlice_l112_355);
  assign when_ArraySlice_l112_355 = (_zz_when_ArraySlice_l112_355 != 6'h0);
  assign when_ArraySlice_l113_355 = (7'h40 <= _zz_when_ArraySlice_l113_355);
  always @(*) begin
    if(when_ArraySlice_l112_355) begin
      if(when_ArraySlice_l113_355) begin
        _zz_when_ArraySlice_l173_355 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_355 = (_zz__zz_when_ArraySlice_l173_355 - _zz__zz_when_ArraySlice_l173_355_3);
      end
    end else begin
      if(when_ArraySlice_l118_355) begin
        _zz_when_ArraySlice_l173_355 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_355 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_355 = (_zz_when_ArraySlice_l118_355 <= wReg);
  assign when_ArraySlice_l173_355 = (_zz_when_ArraySlice_l173_355_1 <= _zz_when_ArraySlice_l173_355_3);
  assign when_ArraySlice_l165_356 = (_zz_when_ArraySlice_l165_356 <= selectWriteFifo);
  assign when_ArraySlice_l166_356 = (_zz_when_ArraySlice_l166_356 <= _zz_when_ArraySlice_l166_356_1);
  assign _zz_when_ArraySlice_l112_356 = (wReg % _zz__zz_when_ArraySlice_l112_356);
  assign when_ArraySlice_l112_356 = (_zz_when_ArraySlice_l112_356 != 6'h0);
  assign when_ArraySlice_l113_356 = (7'h40 <= _zz_when_ArraySlice_l113_356);
  always @(*) begin
    if(when_ArraySlice_l112_356) begin
      if(when_ArraySlice_l113_356) begin
        _zz_when_ArraySlice_l173_356 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_356 = (_zz__zz_when_ArraySlice_l173_356 - _zz__zz_when_ArraySlice_l173_356_3);
      end
    end else begin
      if(when_ArraySlice_l118_356) begin
        _zz_when_ArraySlice_l173_356 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_356 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_356 = (_zz_when_ArraySlice_l118_356 <= wReg);
  assign when_ArraySlice_l173_356 = (_zz_when_ArraySlice_l173_356_1 <= _zz_when_ArraySlice_l173_356_3);
  assign when_ArraySlice_l165_357 = (_zz_when_ArraySlice_l165_357 <= selectWriteFifo);
  assign when_ArraySlice_l166_357 = (_zz_when_ArraySlice_l166_357 <= _zz_when_ArraySlice_l166_357_2);
  assign _zz_when_ArraySlice_l112_357 = (wReg % _zz__zz_when_ArraySlice_l112_357);
  assign when_ArraySlice_l112_357 = (_zz_when_ArraySlice_l112_357 != 6'h0);
  assign when_ArraySlice_l113_357 = (7'h40 <= _zz_when_ArraySlice_l113_357);
  always @(*) begin
    if(when_ArraySlice_l112_357) begin
      if(when_ArraySlice_l113_357) begin
        _zz_when_ArraySlice_l173_357 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_357 = (_zz__zz_when_ArraySlice_l173_357 - _zz__zz_when_ArraySlice_l173_357_3);
      end
    end else begin
      if(when_ArraySlice_l118_357) begin
        _zz_when_ArraySlice_l173_357 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_357 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_357 = (_zz_when_ArraySlice_l118_357 <= wReg);
  assign when_ArraySlice_l173_357 = (_zz_when_ArraySlice_l173_357_1 <= _zz_when_ArraySlice_l173_357_3);
  assign when_ArraySlice_l165_358 = (_zz_when_ArraySlice_l165_358 <= selectWriteFifo);
  assign when_ArraySlice_l166_358 = (_zz_when_ArraySlice_l166_358 <= _zz_when_ArraySlice_l166_358_2);
  assign _zz_when_ArraySlice_l112_358 = (wReg % _zz__zz_when_ArraySlice_l112_358);
  assign when_ArraySlice_l112_358 = (_zz_when_ArraySlice_l112_358 != 6'h0);
  assign when_ArraySlice_l113_358 = (7'h40 <= _zz_when_ArraySlice_l113_358);
  always @(*) begin
    if(when_ArraySlice_l112_358) begin
      if(when_ArraySlice_l113_358) begin
        _zz_when_ArraySlice_l173_358 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_358 = (_zz__zz_when_ArraySlice_l173_358 - _zz__zz_when_ArraySlice_l173_358_3);
      end
    end else begin
      if(when_ArraySlice_l118_358) begin
        _zz_when_ArraySlice_l173_358 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_358 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_358 = (_zz_when_ArraySlice_l118_358 <= wReg);
  assign when_ArraySlice_l173_358 = (_zz_when_ArraySlice_l173_358_1 <= _zz_when_ArraySlice_l173_358_3);
  assign when_ArraySlice_l165_359 = (_zz_when_ArraySlice_l165_359 <= selectWriteFifo);
  assign when_ArraySlice_l166_359 = (_zz_when_ArraySlice_l166_359 <= _zz_when_ArraySlice_l166_359_2);
  assign _zz_when_ArraySlice_l112_359 = (wReg % _zz__zz_when_ArraySlice_l112_359);
  assign when_ArraySlice_l112_359 = (_zz_when_ArraySlice_l112_359 != 6'h0);
  assign when_ArraySlice_l113_359 = (7'h40 <= _zz_when_ArraySlice_l113_359);
  always @(*) begin
    if(when_ArraySlice_l112_359) begin
      if(when_ArraySlice_l113_359) begin
        _zz_when_ArraySlice_l173_359 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_359 = (_zz__zz_when_ArraySlice_l173_359 - _zz__zz_when_ArraySlice_l173_359_3);
      end
    end else begin
      if(when_ArraySlice_l118_359) begin
        _zz_when_ArraySlice_l173_359 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_359 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_359 = (_zz_when_ArraySlice_l118_359 <= wReg);
  assign when_ArraySlice_l173_359 = (_zz_when_ArraySlice_l173_359_1 <= _zz_when_ArraySlice_l173_359_3);
  assign when_ArraySlice_l265_6 = (! ((((((_zz_when_ArraySlice_l265_6 && _zz_when_ArraySlice_l265_6_1) && (holdReadOp_4 == _zz_when_ArraySlice_l265_6_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l265_6_3 && _zz_when_ArraySlice_l265_6_4) && (debug_4_44 == _zz_when_ArraySlice_l265_6_5)) && (debug_5_44 == 1'b1)) && (debug_6_44 == 1'b1)) && (debug_7_44 == 1'b1))));
  assign when_ArraySlice_l268_6 = (wReg <= _zz_when_ArraySlice_l268_6_1);
  assign when_ArraySlice_l272_6 = (_zz_when_ArraySlice_l272_6 == 13'h0);
  assign when_ArraySlice_l276_6 = (_zz_when_ArraySlice_l276_6 == 7'h0);
  assign outputStreamArrayData_6_fire_9 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l277_6 = ((handshakeTimes_6_value == _zz_when_ArraySlice_l277_6) && outputStreamArrayData_6_fire_9);
  assign _zz_when_ArraySlice_l94_43 = (hReg % _zz__zz_when_ArraySlice_l94_43);
  assign when_ArraySlice_l94_43 = (_zz_when_ArraySlice_l94_43 != 6'h0);
  assign when_ArraySlice_l95_43 = (7'h40 <= _zz_when_ArraySlice_l95_43);
  always @(*) begin
    if(when_ArraySlice_l94_43) begin
      if(when_ArraySlice_l95_43) begin
        _zz_when_ArraySlice_l279_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_6 = (_zz__zz_when_ArraySlice_l279_6 - _zz__zz_when_ArraySlice_l279_6_3);
      end
    end else begin
      if(when_ArraySlice_l99_43) begin
        _zz_when_ArraySlice_l279_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_6 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_43 = (_zz_when_ArraySlice_l99_43 <= hReg);
  assign when_ArraySlice_l279_6 = (_zz_when_ArraySlice_l279_6_1 < _zz_when_ArraySlice_l279_6_4);
  always @(*) begin
    debug_0_45 = 1'b0;
    if(when_ArraySlice_l165_360) begin
      if(when_ArraySlice_l166_360) begin
        debug_0_45 = 1'b1;
      end else begin
        debug_0_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_360) begin
        debug_0_45 = 1'b1;
      end else begin
        debug_0_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_45 = 1'b0;
    if(when_ArraySlice_l165_361) begin
      if(when_ArraySlice_l166_361) begin
        debug_1_45 = 1'b1;
      end else begin
        debug_1_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_361) begin
        debug_1_45 = 1'b1;
      end else begin
        debug_1_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_45 = 1'b0;
    if(when_ArraySlice_l165_362) begin
      if(when_ArraySlice_l166_362) begin
        debug_2_45 = 1'b1;
      end else begin
        debug_2_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_362) begin
        debug_2_45 = 1'b1;
      end else begin
        debug_2_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_45 = 1'b0;
    if(when_ArraySlice_l165_363) begin
      if(when_ArraySlice_l166_363) begin
        debug_3_45 = 1'b1;
      end else begin
        debug_3_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_363) begin
        debug_3_45 = 1'b1;
      end else begin
        debug_3_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_45 = 1'b0;
    if(when_ArraySlice_l165_364) begin
      if(when_ArraySlice_l166_364) begin
        debug_4_45 = 1'b1;
      end else begin
        debug_4_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_364) begin
        debug_4_45 = 1'b1;
      end else begin
        debug_4_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_45 = 1'b0;
    if(when_ArraySlice_l165_365) begin
      if(when_ArraySlice_l166_365) begin
        debug_5_45 = 1'b1;
      end else begin
        debug_5_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_365) begin
        debug_5_45 = 1'b1;
      end else begin
        debug_5_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_45 = 1'b0;
    if(when_ArraySlice_l165_366) begin
      if(when_ArraySlice_l166_366) begin
        debug_6_45 = 1'b1;
      end else begin
        debug_6_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_366) begin
        debug_6_45 = 1'b1;
      end else begin
        debug_6_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_45 = 1'b0;
    if(when_ArraySlice_l165_367) begin
      if(when_ArraySlice_l166_367) begin
        debug_7_45 = 1'b1;
      end else begin
        debug_7_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_367) begin
        debug_7_45 = 1'b1;
      end else begin
        debug_7_45 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_360 = (_zz_when_ArraySlice_l165_360 <= selectWriteFifo);
  assign when_ArraySlice_l166_360 = (_zz_when_ArraySlice_l166_360 <= _zz_when_ArraySlice_l166_360_1);
  assign _zz_when_ArraySlice_l112_360 = (wReg % _zz__zz_when_ArraySlice_l112_360);
  assign when_ArraySlice_l112_360 = (_zz_when_ArraySlice_l112_360 != 6'h0);
  assign when_ArraySlice_l113_360 = (7'h40 <= _zz_when_ArraySlice_l113_360);
  always @(*) begin
    if(when_ArraySlice_l112_360) begin
      if(when_ArraySlice_l113_360) begin
        _zz_when_ArraySlice_l173_360 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_360 = (_zz__zz_when_ArraySlice_l173_360 - _zz__zz_when_ArraySlice_l173_360_3);
      end
    end else begin
      if(when_ArraySlice_l118_360) begin
        _zz_when_ArraySlice_l173_360 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_360 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_360 = (_zz_when_ArraySlice_l118_360 <= wReg);
  assign when_ArraySlice_l173_360 = (_zz_when_ArraySlice_l173_360_1 <= _zz_when_ArraySlice_l173_360_2);
  assign when_ArraySlice_l165_361 = (_zz_when_ArraySlice_l165_361 <= selectWriteFifo);
  assign when_ArraySlice_l166_361 = (_zz_when_ArraySlice_l166_361 <= _zz_when_ArraySlice_l166_361_1);
  assign _zz_when_ArraySlice_l112_361 = (wReg % _zz__zz_when_ArraySlice_l112_361);
  assign when_ArraySlice_l112_361 = (_zz_when_ArraySlice_l112_361 != 6'h0);
  assign when_ArraySlice_l113_361 = (7'h40 <= _zz_when_ArraySlice_l113_361);
  always @(*) begin
    if(when_ArraySlice_l112_361) begin
      if(when_ArraySlice_l113_361) begin
        _zz_when_ArraySlice_l173_361 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_361 = (_zz__zz_when_ArraySlice_l173_361 - _zz__zz_when_ArraySlice_l173_361_3);
      end
    end else begin
      if(when_ArraySlice_l118_361) begin
        _zz_when_ArraySlice_l173_361 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_361 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_361 = (_zz_when_ArraySlice_l118_361 <= wReg);
  assign when_ArraySlice_l173_361 = (_zz_when_ArraySlice_l173_361_1 <= _zz_when_ArraySlice_l173_361_3);
  assign when_ArraySlice_l165_362 = (_zz_when_ArraySlice_l165_362 <= selectWriteFifo);
  assign when_ArraySlice_l166_362 = (_zz_when_ArraySlice_l166_362 <= _zz_when_ArraySlice_l166_362_1);
  assign _zz_when_ArraySlice_l112_362 = (wReg % _zz__zz_when_ArraySlice_l112_362);
  assign when_ArraySlice_l112_362 = (_zz_when_ArraySlice_l112_362 != 6'h0);
  assign when_ArraySlice_l113_362 = (7'h40 <= _zz_when_ArraySlice_l113_362);
  always @(*) begin
    if(when_ArraySlice_l112_362) begin
      if(when_ArraySlice_l113_362) begin
        _zz_when_ArraySlice_l173_362 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_362 = (_zz__zz_when_ArraySlice_l173_362 - _zz__zz_when_ArraySlice_l173_362_3);
      end
    end else begin
      if(when_ArraySlice_l118_362) begin
        _zz_when_ArraySlice_l173_362 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_362 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_362 = (_zz_when_ArraySlice_l118_362 <= wReg);
  assign when_ArraySlice_l173_362 = (_zz_when_ArraySlice_l173_362_1 <= _zz_when_ArraySlice_l173_362_3);
  assign when_ArraySlice_l165_363 = (_zz_when_ArraySlice_l165_363 <= selectWriteFifo);
  assign when_ArraySlice_l166_363 = (_zz_when_ArraySlice_l166_363 <= _zz_when_ArraySlice_l166_363_1);
  assign _zz_when_ArraySlice_l112_363 = (wReg % _zz__zz_when_ArraySlice_l112_363);
  assign when_ArraySlice_l112_363 = (_zz_when_ArraySlice_l112_363 != 6'h0);
  assign when_ArraySlice_l113_363 = (7'h40 <= _zz_when_ArraySlice_l113_363);
  always @(*) begin
    if(when_ArraySlice_l112_363) begin
      if(when_ArraySlice_l113_363) begin
        _zz_when_ArraySlice_l173_363 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_363 = (_zz__zz_when_ArraySlice_l173_363 - _zz__zz_when_ArraySlice_l173_363_3);
      end
    end else begin
      if(when_ArraySlice_l118_363) begin
        _zz_when_ArraySlice_l173_363 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_363 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_363 = (_zz_when_ArraySlice_l118_363 <= wReg);
  assign when_ArraySlice_l173_363 = (_zz_when_ArraySlice_l173_363_1 <= _zz_when_ArraySlice_l173_363_3);
  assign when_ArraySlice_l165_364 = (_zz_when_ArraySlice_l165_364 <= selectWriteFifo);
  assign when_ArraySlice_l166_364 = (_zz_when_ArraySlice_l166_364 <= _zz_when_ArraySlice_l166_364_1);
  assign _zz_when_ArraySlice_l112_364 = (wReg % _zz__zz_when_ArraySlice_l112_364);
  assign when_ArraySlice_l112_364 = (_zz_when_ArraySlice_l112_364 != 6'h0);
  assign when_ArraySlice_l113_364 = (7'h40 <= _zz_when_ArraySlice_l113_364);
  always @(*) begin
    if(when_ArraySlice_l112_364) begin
      if(when_ArraySlice_l113_364) begin
        _zz_when_ArraySlice_l173_364 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_364 = (_zz__zz_when_ArraySlice_l173_364 - _zz__zz_when_ArraySlice_l173_364_3);
      end
    end else begin
      if(when_ArraySlice_l118_364) begin
        _zz_when_ArraySlice_l173_364 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_364 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_364 = (_zz_when_ArraySlice_l118_364 <= wReg);
  assign when_ArraySlice_l173_364 = (_zz_when_ArraySlice_l173_364_1 <= _zz_when_ArraySlice_l173_364_3);
  assign when_ArraySlice_l165_365 = (_zz_when_ArraySlice_l165_365 <= selectWriteFifo);
  assign when_ArraySlice_l166_365 = (_zz_when_ArraySlice_l166_365 <= _zz_when_ArraySlice_l166_365_2);
  assign _zz_when_ArraySlice_l112_365 = (wReg % _zz__zz_when_ArraySlice_l112_365);
  assign when_ArraySlice_l112_365 = (_zz_when_ArraySlice_l112_365 != 6'h0);
  assign when_ArraySlice_l113_365 = (7'h40 <= _zz_when_ArraySlice_l113_365);
  always @(*) begin
    if(when_ArraySlice_l112_365) begin
      if(when_ArraySlice_l113_365) begin
        _zz_when_ArraySlice_l173_365 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_365 = (_zz__zz_when_ArraySlice_l173_365 - _zz__zz_when_ArraySlice_l173_365_3);
      end
    end else begin
      if(when_ArraySlice_l118_365) begin
        _zz_when_ArraySlice_l173_365 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_365 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_365 = (_zz_when_ArraySlice_l118_365 <= wReg);
  assign when_ArraySlice_l173_365 = (_zz_when_ArraySlice_l173_365_1 <= _zz_when_ArraySlice_l173_365_3);
  assign when_ArraySlice_l165_366 = (_zz_when_ArraySlice_l165_366 <= selectWriteFifo);
  assign when_ArraySlice_l166_366 = (_zz_when_ArraySlice_l166_366 <= _zz_when_ArraySlice_l166_366_2);
  assign _zz_when_ArraySlice_l112_366 = (wReg % _zz__zz_when_ArraySlice_l112_366);
  assign when_ArraySlice_l112_366 = (_zz_when_ArraySlice_l112_366 != 6'h0);
  assign when_ArraySlice_l113_366 = (7'h40 <= _zz_when_ArraySlice_l113_366);
  always @(*) begin
    if(when_ArraySlice_l112_366) begin
      if(when_ArraySlice_l113_366) begin
        _zz_when_ArraySlice_l173_366 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_366 = (_zz__zz_when_ArraySlice_l173_366 - _zz__zz_when_ArraySlice_l173_366_3);
      end
    end else begin
      if(when_ArraySlice_l118_366) begin
        _zz_when_ArraySlice_l173_366 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_366 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_366 = (_zz_when_ArraySlice_l118_366 <= wReg);
  assign when_ArraySlice_l173_366 = (_zz_when_ArraySlice_l173_366_1 <= _zz_when_ArraySlice_l173_366_3);
  assign when_ArraySlice_l165_367 = (_zz_when_ArraySlice_l165_367 <= selectWriteFifo);
  assign when_ArraySlice_l166_367 = (_zz_when_ArraySlice_l166_367 <= _zz_when_ArraySlice_l166_367_2);
  assign _zz_when_ArraySlice_l112_367 = (wReg % _zz__zz_when_ArraySlice_l112_367);
  assign when_ArraySlice_l112_367 = (_zz_when_ArraySlice_l112_367 != 6'h0);
  assign when_ArraySlice_l113_367 = (7'h40 <= _zz_when_ArraySlice_l113_367);
  always @(*) begin
    if(when_ArraySlice_l112_367) begin
      if(when_ArraySlice_l113_367) begin
        _zz_when_ArraySlice_l173_367 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_367 = (_zz__zz_when_ArraySlice_l173_367 - _zz__zz_when_ArraySlice_l173_367_3);
      end
    end else begin
      if(when_ArraySlice_l118_367) begin
        _zz_when_ArraySlice_l173_367 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_367 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_367 = (_zz_when_ArraySlice_l118_367 <= wReg);
  assign when_ArraySlice_l173_367 = (_zz_when_ArraySlice_l173_367_1 <= _zz_when_ArraySlice_l173_367_3);
  assign when_ArraySlice_l285_6 = (! ((((((_zz_when_ArraySlice_l285_6 && _zz_when_ArraySlice_l285_6_1) && (holdReadOp_4 == _zz_when_ArraySlice_l285_6_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l285_6_3 && _zz_when_ArraySlice_l285_6_4) && (debug_4_45 == _zz_when_ArraySlice_l285_6_5)) && (debug_5_45 == 1'b1)) && (debug_6_45 == 1'b1)) && (debug_7_45 == 1'b1))));
  assign when_ArraySlice_l288_6 = (wReg <= _zz_when_ArraySlice_l288_6_1);
  assign outputStreamArrayData_6_fire_10 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l292_6 = ((_zz_when_ArraySlice_l292_6 == 13'h0) && outputStreamArrayData_6_fire_10);
  assign outputStreamArrayData_6_fire_11 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l303_6 = ((handshakeTimes_6_value == _zz_when_ArraySlice_l303_6) && outputStreamArrayData_6_fire_11);
  assign _zz_when_ArraySlice_l94_44 = (hReg % _zz__zz_when_ArraySlice_l94_44);
  assign when_ArraySlice_l94_44 = (_zz_when_ArraySlice_l94_44 != 6'h0);
  assign when_ArraySlice_l95_44 = (7'h40 <= _zz_when_ArraySlice_l95_44);
  always @(*) begin
    if(when_ArraySlice_l94_44) begin
      if(when_ArraySlice_l95_44) begin
        _zz_when_ArraySlice_l304_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_6 = (_zz__zz_when_ArraySlice_l304_6 - _zz__zz_when_ArraySlice_l304_6_3);
      end
    end else begin
      if(when_ArraySlice_l99_44) begin
        _zz_when_ArraySlice_l304_6 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_6 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_44 = (_zz_when_ArraySlice_l99_44 <= hReg);
  assign when_ArraySlice_l304_6 = (_zz_when_ArraySlice_l304_6_1 < _zz_when_ArraySlice_l304_6_4);
  always @(*) begin
    debug_0_46 = 1'b0;
    if(when_ArraySlice_l165_368) begin
      if(when_ArraySlice_l166_368) begin
        debug_0_46 = 1'b1;
      end else begin
        debug_0_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_368) begin
        debug_0_46 = 1'b1;
      end else begin
        debug_0_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_46 = 1'b0;
    if(when_ArraySlice_l165_369) begin
      if(when_ArraySlice_l166_369) begin
        debug_1_46 = 1'b1;
      end else begin
        debug_1_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_369) begin
        debug_1_46 = 1'b1;
      end else begin
        debug_1_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_46 = 1'b0;
    if(when_ArraySlice_l165_370) begin
      if(when_ArraySlice_l166_370) begin
        debug_2_46 = 1'b1;
      end else begin
        debug_2_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_370) begin
        debug_2_46 = 1'b1;
      end else begin
        debug_2_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_46 = 1'b0;
    if(when_ArraySlice_l165_371) begin
      if(when_ArraySlice_l166_371) begin
        debug_3_46 = 1'b1;
      end else begin
        debug_3_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_371) begin
        debug_3_46 = 1'b1;
      end else begin
        debug_3_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_46 = 1'b0;
    if(when_ArraySlice_l165_372) begin
      if(when_ArraySlice_l166_372) begin
        debug_4_46 = 1'b1;
      end else begin
        debug_4_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_372) begin
        debug_4_46 = 1'b1;
      end else begin
        debug_4_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_46 = 1'b0;
    if(when_ArraySlice_l165_373) begin
      if(when_ArraySlice_l166_373) begin
        debug_5_46 = 1'b1;
      end else begin
        debug_5_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_373) begin
        debug_5_46 = 1'b1;
      end else begin
        debug_5_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_46 = 1'b0;
    if(when_ArraySlice_l165_374) begin
      if(when_ArraySlice_l166_374) begin
        debug_6_46 = 1'b1;
      end else begin
        debug_6_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_374) begin
        debug_6_46 = 1'b1;
      end else begin
        debug_6_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_46 = 1'b0;
    if(when_ArraySlice_l165_375) begin
      if(when_ArraySlice_l166_375) begin
        debug_7_46 = 1'b1;
      end else begin
        debug_7_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_375) begin
        debug_7_46 = 1'b1;
      end else begin
        debug_7_46 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_368 = (_zz_when_ArraySlice_l165_368 <= selectWriteFifo);
  assign when_ArraySlice_l166_368 = (_zz_when_ArraySlice_l166_368 <= _zz_when_ArraySlice_l166_368_1);
  assign _zz_when_ArraySlice_l112_368 = (wReg % _zz__zz_when_ArraySlice_l112_368);
  assign when_ArraySlice_l112_368 = (_zz_when_ArraySlice_l112_368 != 6'h0);
  assign when_ArraySlice_l113_368 = (7'h40 <= _zz_when_ArraySlice_l113_368);
  always @(*) begin
    if(when_ArraySlice_l112_368) begin
      if(when_ArraySlice_l113_368) begin
        _zz_when_ArraySlice_l173_368 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_368 = (_zz__zz_when_ArraySlice_l173_368 - _zz__zz_when_ArraySlice_l173_368_3);
      end
    end else begin
      if(when_ArraySlice_l118_368) begin
        _zz_when_ArraySlice_l173_368 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_368 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_368 = (_zz_when_ArraySlice_l118_368 <= wReg);
  assign when_ArraySlice_l173_368 = (_zz_when_ArraySlice_l173_368_1 <= _zz_when_ArraySlice_l173_368_2);
  assign when_ArraySlice_l165_369 = (_zz_when_ArraySlice_l165_369 <= selectWriteFifo);
  assign when_ArraySlice_l166_369 = (_zz_when_ArraySlice_l166_369 <= _zz_when_ArraySlice_l166_369_1);
  assign _zz_when_ArraySlice_l112_369 = (wReg % _zz__zz_when_ArraySlice_l112_369);
  assign when_ArraySlice_l112_369 = (_zz_when_ArraySlice_l112_369 != 6'h0);
  assign when_ArraySlice_l113_369 = (7'h40 <= _zz_when_ArraySlice_l113_369);
  always @(*) begin
    if(when_ArraySlice_l112_369) begin
      if(when_ArraySlice_l113_369) begin
        _zz_when_ArraySlice_l173_369 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_369 = (_zz__zz_when_ArraySlice_l173_369 - _zz__zz_when_ArraySlice_l173_369_3);
      end
    end else begin
      if(when_ArraySlice_l118_369) begin
        _zz_when_ArraySlice_l173_369 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_369 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_369 = (_zz_when_ArraySlice_l118_369 <= wReg);
  assign when_ArraySlice_l173_369 = (_zz_when_ArraySlice_l173_369_1 <= _zz_when_ArraySlice_l173_369_3);
  assign when_ArraySlice_l165_370 = (_zz_when_ArraySlice_l165_370 <= selectWriteFifo);
  assign when_ArraySlice_l166_370 = (_zz_when_ArraySlice_l166_370 <= _zz_when_ArraySlice_l166_370_1);
  assign _zz_when_ArraySlice_l112_370 = (wReg % _zz__zz_when_ArraySlice_l112_370);
  assign when_ArraySlice_l112_370 = (_zz_when_ArraySlice_l112_370 != 6'h0);
  assign when_ArraySlice_l113_370 = (7'h40 <= _zz_when_ArraySlice_l113_370);
  always @(*) begin
    if(when_ArraySlice_l112_370) begin
      if(when_ArraySlice_l113_370) begin
        _zz_when_ArraySlice_l173_370 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_370 = (_zz__zz_when_ArraySlice_l173_370 - _zz__zz_when_ArraySlice_l173_370_3);
      end
    end else begin
      if(when_ArraySlice_l118_370) begin
        _zz_when_ArraySlice_l173_370 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_370 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_370 = (_zz_when_ArraySlice_l118_370 <= wReg);
  assign when_ArraySlice_l173_370 = (_zz_when_ArraySlice_l173_370_1 <= _zz_when_ArraySlice_l173_370_3);
  assign when_ArraySlice_l165_371 = (_zz_when_ArraySlice_l165_371 <= selectWriteFifo);
  assign when_ArraySlice_l166_371 = (_zz_when_ArraySlice_l166_371 <= _zz_when_ArraySlice_l166_371_1);
  assign _zz_when_ArraySlice_l112_371 = (wReg % _zz__zz_when_ArraySlice_l112_371);
  assign when_ArraySlice_l112_371 = (_zz_when_ArraySlice_l112_371 != 6'h0);
  assign when_ArraySlice_l113_371 = (7'h40 <= _zz_when_ArraySlice_l113_371);
  always @(*) begin
    if(when_ArraySlice_l112_371) begin
      if(when_ArraySlice_l113_371) begin
        _zz_when_ArraySlice_l173_371 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_371 = (_zz__zz_when_ArraySlice_l173_371 - _zz__zz_when_ArraySlice_l173_371_3);
      end
    end else begin
      if(when_ArraySlice_l118_371) begin
        _zz_when_ArraySlice_l173_371 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_371 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_371 = (_zz_when_ArraySlice_l118_371 <= wReg);
  assign when_ArraySlice_l173_371 = (_zz_when_ArraySlice_l173_371_1 <= _zz_when_ArraySlice_l173_371_3);
  assign when_ArraySlice_l165_372 = (_zz_when_ArraySlice_l165_372 <= selectWriteFifo);
  assign when_ArraySlice_l166_372 = (_zz_when_ArraySlice_l166_372 <= _zz_when_ArraySlice_l166_372_1);
  assign _zz_when_ArraySlice_l112_372 = (wReg % _zz__zz_when_ArraySlice_l112_372);
  assign when_ArraySlice_l112_372 = (_zz_when_ArraySlice_l112_372 != 6'h0);
  assign when_ArraySlice_l113_372 = (7'h40 <= _zz_when_ArraySlice_l113_372);
  always @(*) begin
    if(when_ArraySlice_l112_372) begin
      if(when_ArraySlice_l113_372) begin
        _zz_when_ArraySlice_l173_372 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_372 = (_zz__zz_when_ArraySlice_l173_372 - _zz__zz_when_ArraySlice_l173_372_3);
      end
    end else begin
      if(when_ArraySlice_l118_372) begin
        _zz_when_ArraySlice_l173_372 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_372 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_372 = (_zz_when_ArraySlice_l118_372 <= wReg);
  assign when_ArraySlice_l173_372 = (_zz_when_ArraySlice_l173_372_1 <= _zz_when_ArraySlice_l173_372_3);
  assign when_ArraySlice_l165_373 = (_zz_when_ArraySlice_l165_373 <= selectWriteFifo);
  assign when_ArraySlice_l166_373 = (_zz_when_ArraySlice_l166_373 <= _zz_when_ArraySlice_l166_373_2);
  assign _zz_when_ArraySlice_l112_373 = (wReg % _zz__zz_when_ArraySlice_l112_373);
  assign when_ArraySlice_l112_373 = (_zz_when_ArraySlice_l112_373 != 6'h0);
  assign when_ArraySlice_l113_373 = (7'h40 <= _zz_when_ArraySlice_l113_373);
  always @(*) begin
    if(when_ArraySlice_l112_373) begin
      if(when_ArraySlice_l113_373) begin
        _zz_when_ArraySlice_l173_373 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_373 = (_zz__zz_when_ArraySlice_l173_373 - _zz__zz_when_ArraySlice_l173_373_3);
      end
    end else begin
      if(when_ArraySlice_l118_373) begin
        _zz_when_ArraySlice_l173_373 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_373 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_373 = (_zz_when_ArraySlice_l118_373 <= wReg);
  assign when_ArraySlice_l173_373 = (_zz_when_ArraySlice_l173_373_1 <= _zz_when_ArraySlice_l173_373_3);
  assign when_ArraySlice_l165_374 = (_zz_when_ArraySlice_l165_374 <= selectWriteFifo);
  assign when_ArraySlice_l166_374 = (_zz_when_ArraySlice_l166_374 <= _zz_when_ArraySlice_l166_374_2);
  assign _zz_when_ArraySlice_l112_374 = (wReg % _zz__zz_when_ArraySlice_l112_374);
  assign when_ArraySlice_l112_374 = (_zz_when_ArraySlice_l112_374 != 6'h0);
  assign when_ArraySlice_l113_374 = (7'h40 <= _zz_when_ArraySlice_l113_374);
  always @(*) begin
    if(when_ArraySlice_l112_374) begin
      if(when_ArraySlice_l113_374) begin
        _zz_when_ArraySlice_l173_374 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_374 = (_zz__zz_when_ArraySlice_l173_374 - _zz__zz_when_ArraySlice_l173_374_3);
      end
    end else begin
      if(when_ArraySlice_l118_374) begin
        _zz_when_ArraySlice_l173_374 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_374 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_374 = (_zz_when_ArraySlice_l118_374 <= wReg);
  assign when_ArraySlice_l173_374 = (_zz_when_ArraySlice_l173_374_1 <= _zz_when_ArraySlice_l173_374_3);
  assign when_ArraySlice_l165_375 = (_zz_when_ArraySlice_l165_375 <= selectWriteFifo);
  assign when_ArraySlice_l166_375 = (_zz_when_ArraySlice_l166_375 <= _zz_when_ArraySlice_l166_375_2);
  assign _zz_when_ArraySlice_l112_375 = (wReg % _zz__zz_when_ArraySlice_l112_375);
  assign when_ArraySlice_l112_375 = (_zz_when_ArraySlice_l112_375 != 6'h0);
  assign when_ArraySlice_l113_375 = (7'h40 <= _zz_when_ArraySlice_l113_375);
  always @(*) begin
    if(when_ArraySlice_l112_375) begin
      if(when_ArraySlice_l113_375) begin
        _zz_when_ArraySlice_l173_375 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_375 = (_zz__zz_when_ArraySlice_l173_375 - _zz__zz_when_ArraySlice_l173_375_3);
      end
    end else begin
      if(when_ArraySlice_l118_375) begin
        _zz_when_ArraySlice_l173_375 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_375 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_375 = (_zz_when_ArraySlice_l118_375 <= wReg);
  assign when_ArraySlice_l173_375 = (_zz_when_ArraySlice_l173_375_1 <= _zz_when_ArraySlice_l173_375_3);
  assign when_ArraySlice_l311_6 = (! ((((((_zz_when_ArraySlice_l311_6 && _zz_when_ArraySlice_l311_6_1) && (holdReadOp_4 == _zz_when_ArraySlice_l311_6_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l311_6_3 && _zz_when_ArraySlice_l311_6_4) && (debug_4_46 == _zz_when_ArraySlice_l311_6_5)) && (debug_5_46 == 1'b1)) && (debug_6_46 == 1'b1)) && (debug_7_46 == 1'b1))));
  assign outputStreamArrayData_6_fire_12 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l315_6 = ((_zz_when_ArraySlice_l315_6 == 13'h0) && outputStreamArrayData_6_fire_12);
  assign when_ArraySlice_l301_6 = (allowPadding_6 && (wReg <= _zz_when_ArraySlice_l301_6));
  assign outputStreamArrayData_6_fire_13 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l322_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l322_6);
  assign when_ArraySlice_l240_7 = (_zz_when_ArraySlice_l240_7 < wReg);
  assign when_ArraySlice_l241_7 = ((! holdReadOp_7) && (_zz_when_ArraySlice_l241_7 != 7'h0));
  assign _zz_outputStreamArrayData_7_valid_1 = (selectReadFifo_7 + _zz__zz_outputStreamArrayData_7_valid_1);
  assign _zz_18 = ({63'd0,1'b1} <<< _zz_outputStreamArrayData_7_valid_1);
  assign _zz_io_pop_ready_15 = outputStreamArrayData_7_ready;
  assign when_ArraySlice_l246_7 = (! holdReadOp_7);
  assign outputStreamArrayData_7_fire_7 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l247_7 = ((_zz_when_ArraySlice_l247_7 < _zz_when_ArraySlice_l247_7_2) && outputStreamArrayData_7_fire_7);
  assign when_ArraySlice_l248_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l248_7);
  assign when_ArraySlice_l251_7 = (_zz_when_ArraySlice_l251_7 == 13'h0);
  assign outputStreamArrayData_7_fire_8 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l256_7 = ((_zz_when_ArraySlice_l256_7 == _zz_when_ArraySlice_l256_7_3) && outputStreamArrayData_7_fire_8);
  assign when_ArraySlice_l257_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l257_7);
  assign _zz_when_ArraySlice_l94_45 = (hReg % _zz__zz_when_ArraySlice_l94_45);
  assign when_ArraySlice_l94_45 = (_zz_when_ArraySlice_l94_45 != 6'h0);
  assign when_ArraySlice_l95_45 = (7'h40 <= _zz_when_ArraySlice_l95_45);
  always @(*) begin
    if(when_ArraySlice_l94_45) begin
      if(when_ArraySlice_l95_45) begin
        _zz_when_ArraySlice_l259_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_7 = (_zz__zz_when_ArraySlice_l259_7 - _zz__zz_when_ArraySlice_l259_7_3);
      end
    end else begin
      if(when_ArraySlice_l99_45) begin
        _zz_when_ArraySlice_l259_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l259_7 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_45 = (_zz_when_ArraySlice_l99_45 <= hReg);
  assign when_ArraySlice_l259_7 = (_zz_when_ArraySlice_l259_7_1 < _zz_when_ArraySlice_l259_7_4);
  always @(*) begin
    debug_0_47 = 1'b0;
    if(when_ArraySlice_l165_376) begin
      if(when_ArraySlice_l166_376) begin
        debug_0_47 = 1'b1;
      end else begin
        debug_0_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_376) begin
        debug_0_47 = 1'b1;
      end else begin
        debug_0_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_47 = 1'b0;
    if(when_ArraySlice_l165_377) begin
      if(when_ArraySlice_l166_377) begin
        debug_1_47 = 1'b1;
      end else begin
        debug_1_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_377) begin
        debug_1_47 = 1'b1;
      end else begin
        debug_1_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_47 = 1'b0;
    if(when_ArraySlice_l165_378) begin
      if(when_ArraySlice_l166_378) begin
        debug_2_47 = 1'b1;
      end else begin
        debug_2_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_378) begin
        debug_2_47 = 1'b1;
      end else begin
        debug_2_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_47 = 1'b0;
    if(when_ArraySlice_l165_379) begin
      if(when_ArraySlice_l166_379) begin
        debug_3_47 = 1'b1;
      end else begin
        debug_3_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_379) begin
        debug_3_47 = 1'b1;
      end else begin
        debug_3_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_47 = 1'b0;
    if(when_ArraySlice_l165_380) begin
      if(when_ArraySlice_l166_380) begin
        debug_4_47 = 1'b1;
      end else begin
        debug_4_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_380) begin
        debug_4_47 = 1'b1;
      end else begin
        debug_4_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_47 = 1'b0;
    if(when_ArraySlice_l165_381) begin
      if(when_ArraySlice_l166_381) begin
        debug_5_47 = 1'b1;
      end else begin
        debug_5_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_381) begin
        debug_5_47 = 1'b1;
      end else begin
        debug_5_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_47 = 1'b0;
    if(when_ArraySlice_l165_382) begin
      if(when_ArraySlice_l166_382) begin
        debug_6_47 = 1'b1;
      end else begin
        debug_6_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_382) begin
        debug_6_47 = 1'b1;
      end else begin
        debug_6_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_47 = 1'b0;
    if(when_ArraySlice_l165_383) begin
      if(when_ArraySlice_l166_383) begin
        debug_7_47 = 1'b1;
      end else begin
        debug_7_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_383) begin
        debug_7_47 = 1'b1;
      end else begin
        debug_7_47 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_376 = (_zz_when_ArraySlice_l165_376 <= selectWriteFifo);
  assign when_ArraySlice_l166_376 = (_zz_when_ArraySlice_l166_376 <= _zz_when_ArraySlice_l166_376_1);
  assign _zz_when_ArraySlice_l112_376 = (wReg % _zz__zz_when_ArraySlice_l112_376);
  assign when_ArraySlice_l112_376 = (_zz_when_ArraySlice_l112_376 != 6'h0);
  assign when_ArraySlice_l113_376 = (7'h40 <= _zz_when_ArraySlice_l113_376);
  always @(*) begin
    if(when_ArraySlice_l112_376) begin
      if(when_ArraySlice_l113_376) begin
        _zz_when_ArraySlice_l173_376 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_376 = (_zz__zz_when_ArraySlice_l173_376 - _zz__zz_when_ArraySlice_l173_376_3);
      end
    end else begin
      if(when_ArraySlice_l118_376) begin
        _zz_when_ArraySlice_l173_376 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_376 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_376 = (_zz_when_ArraySlice_l118_376 <= wReg);
  assign when_ArraySlice_l173_376 = (_zz_when_ArraySlice_l173_376_1 <= _zz_when_ArraySlice_l173_376_2);
  assign when_ArraySlice_l165_377 = (_zz_when_ArraySlice_l165_377 <= selectWriteFifo);
  assign when_ArraySlice_l166_377 = (_zz_when_ArraySlice_l166_377 <= _zz_when_ArraySlice_l166_377_1);
  assign _zz_when_ArraySlice_l112_377 = (wReg % _zz__zz_when_ArraySlice_l112_377);
  assign when_ArraySlice_l112_377 = (_zz_when_ArraySlice_l112_377 != 6'h0);
  assign when_ArraySlice_l113_377 = (7'h40 <= _zz_when_ArraySlice_l113_377);
  always @(*) begin
    if(when_ArraySlice_l112_377) begin
      if(when_ArraySlice_l113_377) begin
        _zz_when_ArraySlice_l173_377 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_377 = (_zz__zz_when_ArraySlice_l173_377 - _zz__zz_when_ArraySlice_l173_377_3);
      end
    end else begin
      if(when_ArraySlice_l118_377) begin
        _zz_when_ArraySlice_l173_377 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_377 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_377 = (_zz_when_ArraySlice_l118_377 <= wReg);
  assign when_ArraySlice_l173_377 = (_zz_when_ArraySlice_l173_377_1 <= _zz_when_ArraySlice_l173_377_3);
  assign when_ArraySlice_l165_378 = (_zz_when_ArraySlice_l165_378 <= selectWriteFifo);
  assign when_ArraySlice_l166_378 = (_zz_when_ArraySlice_l166_378 <= _zz_when_ArraySlice_l166_378_1);
  assign _zz_when_ArraySlice_l112_378 = (wReg % _zz__zz_when_ArraySlice_l112_378);
  assign when_ArraySlice_l112_378 = (_zz_when_ArraySlice_l112_378 != 6'h0);
  assign when_ArraySlice_l113_378 = (7'h40 <= _zz_when_ArraySlice_l113_378);
  always @(*) begin
    if(when_ArraySlice_l112_378) begin
      if(when_ArraySlice_l113_378) begin
        _zz_when_ArraySlice_l173_378 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_378 = (_zz__zz_when_ArraySlice_l173_378 - _zz__zz_when_ArraySlice_l173_378_3);
      end
    end else begin
      if(when_ArraySlice_l118_378) begin
        _zz_when_ArraySlice_l173_378 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_378 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_378 = (_zz_when_ArraySlice_l118_378 <= wReg);
  assign when_ArraySlice_l173_378 = (_zz_when_ArraySlice_l173_378_1 <= _zz_when_ArraySlice_l173_378_3);
  assign when_ArraySlice_l165_379 = (_zz_when_ArraySlice_l165_379 <= selectWriteFifo);
  assign when_ArraySlice_l166_379 = (_zz_when_ArraySlice_l166_379 <= _zz_when_ArraySlice_l166_379_1);
  assign _zz_when_ArraySlice_l112_379 = (wReg % _zz__zz_when_ArraySlice_l112_379);
  assign when_ArraySlice_l112_379 = (_zz_when_ArraySlice_l112_379 != 6'h0);
  assign when_ArraySlice_l113_379 = (7'h40 <= _zz_when_ArraySlice_l113_379);
  always @(*) begin
    if(when_ArraySlice_l112_379) begin
      if(when_ArraySlice_l113_379) begin
        _zz_when_ArraySlice_l173_379 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_379 = (_zz__zz_when_ArraySlice_l173_379 - _zz__zz_when_ArraySlice_l173_379_3);
      end
    end else begin
      if(when_ArraySlice_l118_379) begin
        _zz_when_ArraySlice_l173_379 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_379 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_379 = (_zz_when_ArraySlice_l118_379 <= wReg);
  assign when_ArraySlice_l173_379 = (_zz_when_ArraySlice_l173_379_1 <= _zz_when_ArraySlice_l173_379_3);
  assign when_ArraySlice_l165_380 = (_zz_when_ArraySlice_l165_380 <= selectWriteFifo);
  assign when_ArraySlice_l166_380 = (_zz_when_ArraySlice_l166_380 <= _zz_when_ArraySlice_l166_380_1);
  assign _zz_when_ArraySlice_l112_380 = (wReg % _zz__zz_when_ArraySlice_l112_380);
  assign when_ArraySlice_l112_380 = (_zz_when_ArraySlice_l112_380 != 6'h0);
  assign when_ArraySlice_l113_380 = (7'h40 <= _zz_when_ArraySlice_l113_380);
  always @(*) begin
    if(when_ArraySlice_l112_380) begin
      if(when_ArraySlice_l113_380) begin
        _zz_when_ArraySlice_l173_380 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_380 = (_zz__zz_when_ArraySlice_l173_380 - _zz__zz_when_ArraySlice_l173_380_3);
      end
    end else begin
      if(when_ArraySlice_l118_380) begin
        _zz_when_ArraySlice_l173_380 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_380 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_380 = (_zz_when_ArraySlice_l118_380 <= wReg);
  assign when_ArraySlice_l173_380 = (_zz_when_ArraySlice_l173_380_1 <= _zz_when_ArraySlice_l173_380_3);
  assign when_ArraySlice_l165_381 = (_zz_when_ArraySlice_l165_381 <= selectWriteFifo);
  assign when_ArraySlice_l166_381 = (_zz_when_ArraySlice_l166_381 <= _zz_when_ArraySlice_l166_381_2);
  assign _zz_when_ArraySlice_l112_381 = (wReg % _zz__zz_when_ArraySlice_l112_381);
  assign when_ArraySlice_l112_381 = (_zz_when_ArraySlice_l112_381 != 6'h0);
  assign when_ArraySlice_l113_381 = (7'h40 <= _zz_when_ArraySlice_l113_381);
  always @(*) begin
    if(when_ArraySlice_l112_381) begin
      if(when_ArraySlice_l113_381) begin
        _zz_when_ArraySlice_l173_381 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_381 = (_zz__zz_when_ArraySlice_l173_381 - _zz__zz_when_ArraySlice_l173_381_3);
      end
    end else begin
      if(when_ArraySlice_l118_381) begin
        _zz_when_ArraySlice_l173_381 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_381 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_381 = (_zz_when_ArraySlice_l118_381 <= wReg);
  assign when_ArraySlice_l173_381 = (_zz_when_ArraySlice_l173_381_1 <= _zz_when_ArraySlice_l173_381_3);
  assign when_ArraySlice_l165_382 = (_zz_when_ArraySlice_l165_382 <= selectWriteFifo);
  assign when_ArraySlice_l166_382 = (_zz_when_ArraySlice_l166_382 <= _zz_when_ArraySlice_l166_382_2);
  assign _zz_when_ArraySlice_l112_382 = (wReg % _zz__zz_when_ArraySlice_l112_382);
  assign when_ArraySlice_l112_382 = (_zz_when_ArraySlice_l112_382 != 6'h0);
  assign when_ArraySlice_l113_382 = (7'h40 <= _zz_when_ArraySlice_l113_382);
  always @(*) begin
    if(when_ArraySlice_l112_382) begin
      if(when_ArraySlice_l113_382) begin
        _zz_when_ArraySlice_l173_382 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_382 = (_zz__zz_when_ArraySlice_l173_382 - _zz__zz_when_ArraySlice_l173_382_3);
      end
    end else begin
      if(when_ArraySlice_l118_382) begin
        _zz_when_ArraySlice_l173_382 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_382 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_382 = (_zz_when_ArraySlice_l118_382 <= wReg);
  assign when_ArraySlice_l173_382 = (_zz_when_ArraySlice_l173_382_1 <= _zz_when_ArraySlice_l173_382_3);
  assign when_ArraySlice_l165_383 = (_zz_when_ArraySlice_l165_383 <= selectWriteFifo);
  assign when_ArraySlice_l166_383 = (_zz_when_ArraySlice_l166_383 <= _zz_when_ArraySlice_l166_383_2);
  assign _zz_when_ArraySlice_l112_383 = (wReg % _zz__zz_when_ArraySlice_l112_383);
  assign when_ArraySlice_l112_383 = (_zz_when_ArraySlice_l112_383 != 6'h0);
  assign when_ArraySlice_l113_383 = (7'h40 <= _zz_when_ArraySlice_l113_383);
  always @(*) begin
    if(when_ArraySlice_l112_383) begin
      if(when_ArraySlice_l113_383) begin
        _zz_when_ArraySlice_l173_383 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_383 = (_zz__zz_when_ArraySlice_l173_383 - _zz__zz_when_ArraySlice_l173_383_3);
      end
    end else begin
      if(when_ArraySlice_l118_383) begin
        _zz_when_ArraySlice_l173_383 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_383 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_383 = (_zz_when_ArraySlice_l118_383 <= wReg);
  assign when_ArraySlice_l173_383 = (_zz_when_ArraySlice_l173_383_1 <= _zz_when_ArraySlice_l173_383_3);
  assign when_ArraySlice_l265_7 = (! ((((((_zz_when_ArraySlice_l265_7 && _zz_when_ArraySlice_l265_7_1) && (holdReadOp_4 == _zz_when_ArraySlice_l265_7_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l265_7_3 && _zz_when_ArraySlice_l265_7_4) && (debug_4_47 == _zz_when_ArraySlice_l265_7_5)) && (debug_5_47 == 1'b1)) && (debug_6_47 == 1'b1)) && (debug_7_47 == 1'b1))));
  assign when_ArraySlice_l268_7 = (wReg <= _zz_when_ArraySlice_l268_7_1);
  assign when_ArraySlice_l272_7 = (_zz_when_ArraySlice_l272_7 == 13'h0);
  assign when_ArraySlice_l276_7 = (_zz_when_ArraySlice_l276_7 == 7'h0);
  assign outputStreamArrayData_7_fire_9 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l277_7 = ((handshakeTimes_7_value == _zz_when_ArraySlice_l277_7) && outputStreamArrayData_7_fire_9);
  assign _zz_when_ArraySlice_l94_46 = (hReg % _zz__zz_when_ArraySlice_l94_46);
  assign when_ArraySlice_l94_46 = (_zz_when_ArraySlice_l94_46 != 6'h0);
  assign when_ArraySlice_l95_46 = (7'h40 <= _zz_when_ArraySlice_l95_46);
  always @(*) begin
    if(when_ArraySlice_l94_46) begin
      if(when_ArraySlice_l95_46) begin
        _zz_when_ArraySlice_l279_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_7 = (_zz__zz_when_ArraySlice_l279_7 - _zz__zz_when_ArraySlice_l279_7_3);
      end
    end else begin
      if(when_ArraySlice_l99_46) begin
        _zz_when_ArraySlice_l279_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l279_7 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_46 = (_zz_when_ArraySlice_l99_46 <= hReg);
  assign when_ArraySlice_l279_7 = (_zz_when_ArraySlice_l279_7_1 < _zz_when_ArraySlice_l279_7_4);
  always @(*) begin
    debug_0_48 = 1'b0;
    if(when_ArraySlice_l165_384) begin
      if(when_ArraySlice_l166_384) begin
        debug_0_48 = 1'b1;
      end else begin
        debug_0_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_384) begin
        debug_0_48 = 1'b1;
      end else begin
        debug_0_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_48 = 1'b0;
    if(when_ArraySlice_l165_385) begin
      if(when_ArraySlice_l166_385) begin
        debug_1_48 = 1'b1;
      end else begin
        debug_1_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_385) begin
        debug_1_48 = 1'b1;
      end else begin
        debug_1_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_48 = 1'b0;
    if(when_ArraySlice_l165_386) begin
      if(when_ArraySlice_l166_386) begin
        debug_2_48 = 1'b1;
      end else begin
        debug_2_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_386) begin
        debug_2_48 = 1'b1;
      end else begin
        debug_2_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_48 = 1'b0;
    if(when_ArraySlice_l165_387) begin
      if(when_ArraySlice_l166_387) begin
        debug_3_48 = 1'b1;
      end else begin
        debug_3_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_387) begin
        debug_3_48 = 1'b1;
      end else begin
        debug_3_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_48 = 1'b0;
    if(when_ArraySlice_l165_388) begin
      if(when_ArraySlice_l166_388) begin
        debug_4_48 = 1'b1;
      end else begin
        debug_4_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_388) begin
        debug_4_48 = 1'b1;
      end else begin
        debug_4_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_48 = 1'b0;
    if(when_ArraySlice_l165_389) begin
      if(when_ArraySlice_l166_389) begin
        debug_5_48 = 1'b1;
      end else begin
        debug_5_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_389) begin
        debug_5_48 = 1'b1;
      end else begin
        debug_5_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_48 = 1'b0;
    if(when_ArraySlice_l165_390) begin
      if(when_ArraySlice_l166_390) begin
        debug_6_48 = 1'b1;
      end else begin
        debug_6_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_390) begin
        debug_6_48 = 1'b1;
      end else begin
        debug_6_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_48 = 1'b0;
    if(when_ArraySlice_l165_391) begin
      if(when_ArraySlice_l166_391) begin
        debug_7_48 = 1'b1;
      end else begin
        debug_7_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_391) begin
        debug_7_48 = 1'b1;
      end else begin
        debug_7_48 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_384 = (_zz_when_ArraySlice_l165_384 <= selectWriteFifo);
  assign when_ArraySlice_l166_384 = (_zz_when_ArraySlice_l166_384 <= _zz_when_ArraySlice_l166_384_1);
  assign _zz_when_ArraySlice_l112_384 = (wReg % _zz__zz_when_ArraySlice_l112_384);
  assign when_ArraySlice_l112_384 = (_zz_when_ArraySlice_l112_384 != 6'h0);
  assign when_ArraySlice_l113_384 = (7'h40 <= _zz_when_ArraySlice_l113_384);
  always @(*) begin
    if(when_ArraySlice_l112_384) begin
      if(when_ArraySlice_l113_384) begin
        _zz_when_ArraySlice_l173_384 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_384 = (_zz__zz_when_ArraySlice_l173_384 - _zz__zz_when_ArraySlice_l173_384_3);
      end
    end else begin
      if(when_ArraySlice_l118_384) begin
        _zz_when_ArraySlice_l173_384 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_384 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_384 = (_zz_when_ArraySlice_l118_384 <= wReg);
  assign when_ArraySlice_l173_384 = (_zz_when_ArraySlice_l173_384_1 <= _zz_when_ArraySlice_l173_384_2);
  assign when_ArraySlice_l165_385 = (_zz_when_ArraySlice_l165_385 <= selectWriteFifo);
  assign when_ArraySlice_l166_385 = (_zz_when_ArraySlice_l166_385 <= _zz_when_ArraySlice_l166_385_1);
  assign _zz_when_ArraySlice_l112_385 = (wReg % _zz__zz_when_ArraySlice_l112_385);
  assign when_ArraySlice_l112_385 = (_zz_when_ArraySlice_l112_385 != 6'h0);
  assign when_ArraySlice_l113_385 = (7'h40 <= _zz_when_ArraySlice_l113_385);
  always @(*) begin
    if(when_ArraySlice_l112_385) begin
      if(when_ArraySlice_l113_385) begin
        _zz_when_ArraySlice_l173_385 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_385 = (_zz__zz_when_ArraySlice_l173_385 - _zz__zz_when_ArraySlice_l173_385_3);
      end
    end else begin
      if(when_ArraySlice_l118_385) begin
        _zz_when_ArraySlice_l173_385 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_385 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_385 = (_zz_when_ArraySlice_l118_385 <= wReg);
  assign when_ArraySlice_l173_385 = (_zz_when_ArraySlice_l173_385_1 <= _zz_when_ArraySlice_l173_385_3);
  assign when_ArraySlice_l165_386 = (_zz_when_ArraySlice_l165_386 <= selectWriteFifo);
  assign when_ArraySlice_l166_386 = (_zz_when_ArraySlice_l166_386 <= _zz_when_ArraySlice_l166_386_1);
  assign _zz_when_ArraySlice_l112_386 = (wReg % _zz__zz_when_ArraySlice_l112_386);
  assign when_ArraySlice_l112_386 = (_zz_when_ArraySlice_l112_386 != 6'h0);
  assign when_ArraySlice_l113_386 = (7'h40 <= _zz_when_ArraySlice_l113_386);
  always @(*) begin
    if(when_ArraySlice_l112_386) begin
      if(when_ArraySlice_l113_386) begin
        _zz_when_ArraySlice_l173_386 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_386 = (_zz__zz_when_ArraySlice_l173_386 - _zz__zz_when_ArraySlice_l173_386_3);
      end
    end else begin
      if(when_ArraySlice_l118_386) begin
        _zz_when_ArraySlice_l173_386 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_386 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_386 = (_zz_when_ArraySlice_l118_386 <= wReg);
  assign when_ArraySlice_l173_386 = (_zz_when_ArraySlice_l173_386_1 <= _zz_when_ArraySlice_l173_386_3);
  assign when_ArraySlice_l165_387 = (_zz_when_ArraySlice_l165_387 <= selectWriteFifo);
  assign when_ArraySlice_l166_387 = (_zz_when_ArraySlice_l166_387 <= _zz_when_ArraySlice_l166_387_1);
  assign _zz_when_ArraySlice_l112_387 = (wReg % _zz__zz_when_ArraySlice_l112_387);
  assign when_ArraySlice_l112_387 = (_zz_when_ArraySlice_l112_387 != 6'h0);
  assign when_ArraySlice_l113_387 = (7'h40 <= _zz_when_ArraySlice_l113_387);
  always @(*) begin
    if(when_ArraySlice_l112_387) begin
      if(when_ArraySlice_l113_387) begin
        _zz_when_ArraySlice_l173_387 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_387 = (_zz__zz_when_ArraySlice_l173_387 - _zz__zz_when_ArraySlice_l173_387_3);
      end
    end else begin
      if(when_ArraySlice_l118_387) begin
        _zz_when_ArraySlice_l173_387 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_387 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_387 = (_zz_when_ArraySlice_l118_387 <= wReg);
  assign when_ArraySlice_l173_387 = (_zz_when_ArraySlice_l173_387_1 <= _zz_when_ArraySlice_l173_387_3);
  assign when_ArraySlice_l165_388 = (_zz_when_ArraySlice_l165_388 <= selectWriteFifo);
  assign when_ArraySlice_l166_388 = (_zz_when_ArraySlice_l166_388 <= _zz_when_ArraySlice_l166_388_1);
  assign _zz_when_ArraySlice_l112_388 = (wReg % _zz__zz_when_ArraySlice_l112_388);
  assign when_ArraySlice_l112_388 = (_zz_when_ArraySlice_l112_388 != 6'h0);
  assign when_ArraySlice_l113_388 = (7'h40 <= _zz_when_ArraySlice_l113_388);
  always @(*) begin
    if(when_ArraySlice_l112_388) begin
      if(when_ArraySlice_l113_388) begin
        _zz_when_ArraySlice_l173_388 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_388 = (_zz__zz_when_ArraySlice_l173_388 - _zz__zz_when_ArraySlice_l173_388_3);
      end
    end else begin
      if(when_ArraySlice_l118_388) begin
        _zz_when_ArraySlice_l173_388 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_388 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_388 = (_zz_when_ArraySlice_l118_388 <= wReg);
  assign when_ArraySlice_l173_388 = (_zz_when_ArraySlice_l173_388_1 <= _zz_when_ArraySlice_l173_388_3);
  assign when_ArraySlice_l165_389 = (_zz_when_ArraySlice_l165_389 <= selectWriteFifo);
  assign when_ArraySlice_l166_389 = (_zz_when_ArraySlice_l166_389 <= _zz_when_ArraySlice_l166_389_2);
  assign _zz_when_ArraySlice_l112_389 = (wReg % _zz__zz_when_ArraySlice_l112_389);
  assign when_ArraySlice_l112_389 = (_zz_when_ArraySlice_l112_389 != 6'h0);
  assign when_ArraySlice_l113_389 = (7'h40 <= _zz_when_ArraySlice_l113_389);
  always @(*) begin
    if(when_ArraySlice_l112_389) begin
      if(when_ArraySlice_l113_389) begin
        _zz_when_ArraySlice_l173_389 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_389 = (_zz__zz_when_ArraySlice_l173_389 - _zz__zz_when_ArraySlice_l173_389_3);
      end
    end else begin
      if(when_ArraySlice_l118_389) begin
        _zz_when_ArraySlice_l173_389 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_389 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_389 = (_zz_when_ArraySlice_l118_389 <= wReg);
  assign when_ArraySlice_l173_389 = (_zz_when_ArraySlice_l173_389_1 <= _zz_when_ArraySlice_l173_389_3);
  assign when_ArraySlice_l165_390 = (_zz_when_ArraySlice_l165_390 <= selectWriteFifo);
  assign when_ArraySlice_l166_390 = (_zz_when_ArraySlice_l166_390 <= _zz_when_ArraySlice_l166_390_2);
  assign _zz_when_ArraySlice_l112_390 = (wReg % _zz__zz_when_ArraySlice_l112_390);
  assign when_ArraySlice_l112_390 = (_zz_when_ArraySlice_l112_390 != 6'h0);
  assign when_ArraySlice_l113_390 = (7'h40 <= _zz_when_ArraySlice_l113_390);
  always @(*) begin
    if(when_ArraySlice_l112_390) begin
      if(when_ArraySlice_l113_390) begin
        _zz_when_ArraySlice_l173_390 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_390 = (_zz__zz_when_ArraySlice_l173_390 - _zz__zz_when_ArraySlice_l173_390_3);
      end
    end else begin
      if(when_ArraySlice_l118_390) begin
        _zz_when_ArraySlice_l173_390 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_390 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_390 = (_zz_when_ArraySlice_l118_390 <= wReg);
  assign when_ArraySlice_l173_390 = (_zz_when_ArraySlice_l173_390_1 <= _zz_when_ArraySlice_l173_390_3);
  assign when_ArraySlice_l165_391 = (_zz_when_ArraySlice_l165_391 <= selectWriteFifo);
  assign when_ArraySlice_l166_391 = (_zz_when_ArraySlice_l166_391 <= _zz_when_ArraySlice_l166_391_2);
  assign _zz_when_ArraySlice_l112_391 = (wReg % _zz__zz_when_ArraySlice_l112_391);
  assign when_ArraySlice_l112_391 = (_zz_when_ArraySlice_l112_391 != 6'h0);
  assign when_ArraySlice_l113_391 = (7'h40 <= _zz_when_ArraySlice_l113_391);
  always @(*) begin
    if(when_ArraySlice_l112_391) begin
      if(when_ArraySlice_l113_391) begin
        _zz_when_ArraySlice_l173_391 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_391 = (_zz__zz_when_ArraySlice_l173_391 - _zz__zz_when_ArraySlice_l173_391_3);
      end
    end else begin
      if(when_ArraySlice_l118_391) begin
        _zz_when_ArraySlice_l173_391 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_391 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_391 = (_zz_when_ArraySlice_l118_391 <= wReg);
  assign when_ArraySlice_l173_391 = (_zz_when_ArraySlice_l173_391_1 <= _zz_when_ArraySlice_l173_391_3);
  assign when_ArraySlice_l285_7 = (! ((((((_zz_when_ArraySlice_l285_7 && _zz_when_ArraySlice_l285_7_1) && (holdReadOp_4 == _zz_when_ArraySlice_l285_7_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l285_7_3 && _zz_when_ArraySlice_l285_7_4) && (debug_4_48 == _zz_when_ArraySlice_l285_7_5)) && (debug_5_48 == 1'b1)) && (debug_6_48 == 1'b1)) && (debug_7_48 == 1'b1))));
  assign when_ArraySlice_l288_7 = (wReg <= _zz_when_ArraySlice_l288_7_1);
  assign outputStreamArrayData_7_fire_10 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l292_7 = ((_zz_when_ArraySlice_l292_7 == 13'h0) && outputStreamArrayData_7_fire_10);
  assign outputStreamArrayData_7_fire_11 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l303_7 = ((handshakeTimes_7_value == _zz_when_ArraySlice_l303_7) && outputStreamArrayData_7_fire_11);
  assign _zz_when_ArraySlice_l94_47 = (hReg % _zz__zz_when_ArraySlice_l94_47);
  assign when_ArraySlice_l94_47 = (_zz_when_ArraySlice_l94_47 != 6'h0);
  assign when_ArraySlice_l95_47 = (7'h40 <= _zz_when_ArraySlice_l95_47);
  always @(*) begin
    if(when_ArraySlice_l94_47) begin
      if(when_ArraySlice_l95_47) begin
        _zz_when_ArraySlice_l304_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_7 = (_zz__zz_when_ArraySlice_l304_7 - _zz__zz_when_ArraySlice_l304_7_3);
      end
    end else begin
      if(when_ArraySlice_l99_47) begin
        _zz_when_ArraySlice_l304_7 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l304_7 = {1'd0, hReg};
      end
    end
  end

  assign when_ArraySlice_l99_47 = (_zz_when_ArraySlice_l99_47 <= hReg);
  assign when_ArraySlice_l304_7 = (_zz_when_ArraySlice_l304_7_1 < _zz_when_ArraySlice_l304_7_4);
  always @(*) begin
    debug_0_49 = 1'b0;
    if(when_ArraySlice_l165_392) begin
      if(when_ArraySlice_l166_392) begin
        debug_0_49 = 1'b1;
      end else begin
        debug_0_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_392) begin
        debug_0_49 = 1'b1;
      end else begin
        debug_0_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_49 = 1'b0;
    if(when_ArraySlice_l165_393) begin
      if(when_ArraySlice_l166_393) begin
        debug_1_49 = 1'b1;
      end else begin
        debug_1_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_393) begin
        debug_1_49 = 1'b1;
      end else begin
        debug_1_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_49 = 1'b0;
    if(when_ArraySlice_l165_394) begin
      if(when_ArraySlice_l166_394) begin
        debug_2_49 = 1'b1;
      end else begin
        debug_2_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_394) begin
        debug_2_49 = 1'b1;
      end else begin
        debug_2_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_49 = 1'b0;
    if(when_ArraySlice_l165_395) begin
      if(when_ArraySlice_l166_395) begin
        debug_3_49 = 1'b1;
      end else begin
        debug_3_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_395) begin
        debug_3_49 = 1'b1;
      end else begin
        debug_3_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_49 = 1'b0;
    if(when_ArraySlice_l165_396) begin
      if(when_ArraySlice_l166_396) begin
        debug_4_49 = 1'b1;
      end else begin
        debug_4_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_396) begin
        debug_4_49 = 1'b1;
      end else begin
        debug_4_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_49 = 1'b0;
    if(when_ArraySlice_l165_397) begin
      if(when_ArraySlice_l166_397) begin
        debug_5_49 = 1'b1;
      end else begin
        debug_5_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_397) begin
        debug_5_49 = 1'b1;
      end else begin
        debug_5_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_49 = 1'b0;
    if(when_ArraySlice_l165_398) begin
      if(when_ArraySlice_l166_398) begin
        debug_6_49 = 1'b1;
      end else begin
        debug_6_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_398) begin
        debug_6_49 = 1'b1;
      end else begin
        debug_6_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_49 = 1'b0;
    if(when_ArraySlice_l165_399) begin
      if(when_ArraySlice_l166_399) begin
        debug_7_49 = 1'b1;
      end else begin
        debug_7_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_399) begin
        debug_7_49 = 1'b1;
      end else begin
        debug_7_49 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_392 = (_zz_when_ArraySlice_l165_392 <= selectWriteFifo);
  assign when_ArraySlice_l166_392 = (_zz_when_ArraySlice_l166_392 <= _zz_when_ArraySlice_l166_392_1);
  assign _zz_when_ArraySlice_l112_392 = (wReg % _zz__zz_when_ArraySlice_l112_392);
  assign when_ArraySlice_l112_392 = (_zz_when_ArraySlice_l112_392 != 6'h0);
  assign when_ArraySlice_l113_392 = (7'h40 <= _zz_when_ArraySlice_l113_392);
  always @(*) begin
    if(when_ArraySlice_l112_392) begin
      if(when_ArraySlice_l113_392) begin
        _zz_when_ArraySlice_l173_392 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_392 = (_zz__zz_when_ArraySlice_l173_392 - _zz__zz_when_ArraySlice_l173_392_3);
      end
    end else begin
      if(when_ArraySlice_l118_392) begin
        _zz_when_ArraySlice_l173_392 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_392 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_392 = (_zz_when_ArraySlice_l118_392 <= wReg);
  assign when_ArraySlice_l173_392 = (_zz_when_ArraySlice_l173_392_1 <= _zz_when_ArraySlice_l173_392_2);
  assign when_ArraySlice_l165_393 = (_zz_when_ArraySlice_l165_393 <= selectWriteFifo);
  assign when_ArraySlice_l166_393 = (_zz_when_ArraySlice_l166_393 <= _zz_when_ArraySlice_l166_393_1);
  assign _zz_when_ArraySlice_l112_393 = (wReg % _zz__zz_when_ArraySlice_l112_393);
  assign when_ArraySlice_l112_393 = (_zz_when_ArraySlice_l112_393 != 6'h0);
  assign when_ArraySlice_l113_393 = (7'h40 <= _zz_when_ArraySlice_l113_393);
  always @(*) begin
    if(when_ArraySlice_l112_393) begin
      if(when_ArraySlice_l113_393) begin
        _zz_when_ArraySlice_l173_393 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_393 = (_zz__zz_when_ArraySlice_l173_393 - _zz__zz_when_ArraySlice_l173_393_3);
      end
    end else begin
      if(when_ArraySlice_l118_393) begin
        _zz_when_ArraySlice_l173_393 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_393 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_393 = (_zz_when_ArraySlice_l118_393 <= wReg);
  assign when_ArraySlice_l173_393 = (_zz_when_ArraySlice_l173_393_1 <= _zz_when_ArraySlice_l173_393_3);
  assign when_ArraySlice_l165_394 = (_zz_when_ArraySlice_l165_394 <= selectWriteFifo);
  assign when_ArraySlice_l166_394 = (_zz_when_ArraySlice_l166_394 <= _zz_when_ArraySlice_l166_394_1);
  assign _zz_when_ArraySlice_l112_394 = (wReg % _zz__zz_when_ArraySlice_l112_394);
  assign when_ArraySlice_l112_394 = (_zz_when_ArraySlice_l112_394 != 6'h0);
  assign when_ArraySlice_l113_394 = (7'h40 <= _zz_when_ArraySlice_l113_394);
  always @(*) begin
    if(when_ArraySlice_l112_394) begin
      if(when_ArraySlice_l113_394) begin
        _zz_when_ArraySlice_l173_394 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_394 = (_zz__zz_when_ArraySlice_l173_394 - _zz__zz_when_ArraySlice_l173_394_3);
      end
    end else begin
      if(when_ArraySlice_l118_394) begin
        _zz_when_ArraySlice_l173_394 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_394 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_394 = (_zz_when_ArraySlice_l118_394 <= wReg);
  assign when_ArraySlice_l173_394 = (_zz_when_ArraySlice_l173_394_1 <= _zz_when_ArraySlice_l173_394_3);
  assign when_ArraySlice_l165_395 = (_zz_when_ArraySlice_l165_395 <= selectWriteFifo);
  assign when_ArraySlice_l166_395 = (_zz_when_ArraySlice_l166_395 <= _zz_when_ArraySlice_l166_395_1);
  assign _zz_when_ArraySlice_l112_395 = (wReg % _zz__zz_when_ArraySlice_l112_395);
  assign when_ArraySlice_l112_395 = (_zz_when_ArraySlice_l112_395 != 6'h0);
  assign when_ArraySlice_l113_395 = (7'h40 <= _zz_when_ArraySlice_l113_395);
  always @(*) begin
    if(when_ArraySlice_l112_395) begin
      if(when_ArraySlice_l113_395) begin
        _zz_when_ArraySlice_l173_395 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_395 = (_zz__zz_when_ArraySlice_l173_395 - _zz__zz_when_ArraySlice_l173_395_3);
      end
    end else begin
      if(when_ArraySlice_l118_395) begin
        _zz_when_ArraySlice_l173_395 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_395 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_395 = (_zz_when_ArraySlice_l118_395 <= wReg);
  assign when_ArraySlice_l173_395 = (_zz_when_ArraySlice_l173_395_1 <= _zz_when_ArraySlice_l173_395_3);
  assign when_ArraySlice_l165_396 = (_zz_when_ArraySlice_l165_396 <= selectWriteFifo);
  assign when_ArraySlice_l166_396 = (_zz_when_ArraySlice_l166_396 <= _zz_when_ArraySlice_l166_396_1);
  assign _zz_when_ArraySlice_l112_396 = (wReg % _zz__zz_when_ArraySlice_l112_396);
  assign when_ArraySlice_l112_396 = (_zz_when_ArraySlice_l112_396 != 6'h0);
  assign when_ArraySlice_l113_396 = (7'h40 <= _zz_when_ArraySlice_l113_396);
  always @(*) begin
    if(when_ArraySlice_l112_396) begin
      if(when_ArraySlice_l113_396) begin
        _zz_when_ArraySlice_l173_396 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_396 = (_zz__zz_when_ArraySlice_l173_396 - _zz__zz_when_ArraySlice_l173_396_3);
      end
    end else begin
      if(when_ArraySlice_l118_396) begin
        _zz_when_ArraySlice_l173_396 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_396 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_396 = (_zz_when_ArraySlice_l118_396 <= wReg);
  assign when_ArraySlice_l173_396 = (_zz_when_ArraySlice_l173_396_1 <= _zz_when_ArraySlice_l173_396_3);
  assign when_ArraySlice_l165_397 = (_zz_when_ArraySlice_l165_397 <= selectWriteFifo);
  assign when_ArraySlice_l166_397 = (_zz_when_ArraySlice_l166_397 <= _zz_when_ArraySlice_l166_397_2);
  assign _zz_when_ArraySlice_l112_397 = (wReg % _zz__zz_when_ArraySlice_l112_397);
  assign when_ArraySlice_l112_397 = (_zz_when_ArraySlice_l112_397 != 6'h0);
  assign when_ArraySlice_l113_397 = (7'h40 <= _zz_when_ArraySlice_l113_397);
  always @(*) begin
    if(when_ArraySlice_l112_397) begin
      if(when_ArraySlice_l113_397) begin
        _zz_when_ArraySlice_l173_397 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_397 = (_zz__zz_when_ArraySlice_l173_397 - _zz__zz_when_ArraySlice_l173_397_3);
      end
    end else begin
      if(when_ArraySlice_l118_397) begin
        _zz_when_ArraySlice_l173_397 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_397 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_397 = (_zz_when_ArraySlice_l118_397 <= wReg);
  assign when_ArraySlice_l173_397 = (_zz_when_ArraySlice_l173_397_1 <= _zz_when_ArraySlice_l173_397_3);
  assign when_ArraySlice_l165_398 = (_zz_when_ArraySlice_l165_398 <= selectWriteFifo);
  assign when_ArraySlice_l166_398 = (_zz_when_ArraySlice_l166_398 <= _zz_when_ArraySlice_l166_398_2);
  assign _zz_when_ArraySlice_l112_398 = (wReg % _zz__zz_when_ArraySlice_l112_398);
  assign when_ArraySlice_l112_398 = (_zz_when_ArraySlice_l112_398 != 6'h0);
  assign when_ArraySlice_l113_398 = (7'h40 <= _zz_when_ArraySlice_l113_398);
  always @(*) begin
    if(when_ArraySlice_l112_398) begin
      if(when_ArraySlice_l113_398) begin
        _zz_when_ArraySlice_l173_398 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_398 = (_zz__zz_when_ArraySlice_l173_398 - _zz__zz_when_ArraySlice_l173_398_3);
      end
    end else begin
      if(when_ArraySlice_l118_398) begin
        _zz_when_ArraySlice_l173_398 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_398 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_398 = (_zz_when_ArraySlice_l118_398 <= wReg);
  assign when_ArraySlice_l173_398 = (_zz_when_ArraySlice_l173_398_1 <= _zz_when_ArraySlice_l173_398_3);
  assign when_ArraySlice_l165_399 = (_zz_when_ArraySlice_l165_399 <= selectWriteFifo);
  assign when_ArraySlice_l166_399 = (_zz_when_ArraySlice_l166_399 <= _zz_when_ArraySlice_l166_399_2);
  assign _zz_when_ArraySlice_l112_399 = (wReg % _zz__zz_when_ArraySlice_l112_399);
  assign when_ArraySlice_l112_399 = (_zz_when_ArraySlice_l112_399 != 6'h0);
  assign when_ArraySlice_l113_399 = (7'h40 <= _zz_when_ArraySlice_l113_399);
  always @(*) begin
    if(when_ArraySlice_l112_399) begin
      if(when_ArraySlice_l113_399) begin
        _zz_when_ArraySlice_l173_399 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_399 = (_zz__zz_when_ArraySlice_l173_399 - _zz__zz_when_ArraySlice_l173_399_3);
      end
    end else begin
      if(when_ArraySlice_l118_399) begin
        _zz_when_ArraySlice_l173_399 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_399 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_399 = (_zz_when_ArraySlice_l118_399 <= wReg);
  assign when_ArraySlice_l173_399 = (_zz_when_ArraySlice_l173_399_1 <= _zz_when_ArraySlice_l173_399_3);
  assign when_ArraySlice_l311_7 = (! ((((((_zz_when_ArraySlice_l311_7 && _zz_when_ArraySlice_l311_7_1) && (holdReadOp_4 == _zz_when_ArraySlice_l311_7_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l311_7_3 && _zz_when_ArraySlice_l311_7_4) && (debug_4_49 == _zz_when_ArraySlice_l311_7_5)) && (debug_5_49 == 1'b1)) && (debug_6_49 == 1'b1)) && (debug_7_49 == 1'b1))));
  assign outputStreamArrayData_7_fire_12 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l315_7 = ((_zz_when_ArraySlice_l315_7 == 13'h0) && outputStreamArrayData_7_fire_12);
  assign when_ArraySlice_l301_7 = (allowPadding_7 && (wReg <= _zz_when_ArraySlice_l301_7));
  assign outputStreamArrayData_7_fire_13 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l322_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l322_7);
  assign when_ArraySlice_l189 = (selectWriteFifo == _zz_when_ArraySlice_l189);
  assign when_ArraySlice_l190 = (writeAround ^ readAround_0);
  always @(*) begin
    if(when_ArraySlice_l189) begin
      if(when_ArraySlice_l190) begin
        _zz_when_ArraySlice_l333 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l333 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l333 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_1 = (selectWriteFifo == _zz_when_ArraySlice_l189_1_1);
  assign when_ArraySlice_l190_1 = (writeAround ^ readAround_1);
  always @(*) begin
    if(when_ArraySlice_l189_1) begin
      if(when_ArraySlice_l190_1) begin
        _zz_when_ArraySlice_l333_1 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l333_1 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l333_1 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_2 = (selectWriteFifo == _zz_when_ArraySlice_l189_2);
  assign when_ArraySlice_l190_2 = (writeAround ^ readAround_2);
  always @(*) begin
    if(when_ArraySlice_l189_2) begin
      if(when_ArraySlice_l190_2) begin
        _zz_when_ArraySlice_l333_2 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l333_2 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l333_2 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_3 = (selectWriteFifo == _zz_when_ArraySlice_l189_3);
  assign when_ArraySlice_l190_3 = (writeAround ^ readAround_3);
  always @(*) begin
    if(when_ArraySlice_l189_3) begin
      if(when_ArraySlice_l190_3) begin
        _zz_when_ArraySlice_l333_3 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l333_3 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l333_3 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_4 = (selectWriteFifo == _zz_when_ArraySlice_l189_4);
  assign when_ArraySlice_l190_4 = (writeAround ^ readAround_4);
  always @(*) begin
    if(when_ArraySlice_l189_4) begin
      if(when_ArraySlice_l190_4) begin
        _zz_when_ArraySlice_l333_4 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l333_4 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l333_4 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_5 = (selectWriteFifo == _zz_when_ArraySlice_l189_5);
  assign when_ArraySlice_l190_5 = (writeAround ^ readAround_5);
  always @(*) begin
    if(when_ArraySlice_l189_5) begin
      if(when_ArraySlice_l190_5) begin
        _zz_when_ArraySlice_l333_5 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l333_5 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l333_5 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_6 = (selectWriteFifo == _zz_when_ArraySlice_l189_6);
  assign when_ArraySlice_l190_6 = (writeAround ^ readAround_6);
  always @(*) begin
    if(when_ArraySlice_l189_6) begin
      if(when_ArraySlice_l190_6) begin
        _zz_when_ArraySlice_l333_6 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l333_6 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l333_6 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_7 = (selectWriteFifo == _zz_when_ArraySlice_l189_7);
  assign when_ArraySlice_l190_7 = (writeAround ^ readAround_7);
  always @(*) begin
    if(when_ArraySlice_l189_7) begin
      if(when_ArraySlice_l190_7) begin
        _zz_when_ArraySlice_l333_7 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l333_7 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l333_7 = 1'b0;
    end
  end

  assign when_ArraySlice_l333 = (! ((((((((_zz_when_ArraySlice_l333 != _zz_when_ArraySlice_l333_8) || (_zz_when_ArraySlice_l333_1 != _zz_when_ArraySlice_l333_9)) || (_zz_when_ArraySlice_l333_2 != 1'b0)) || (_zz_when_ArraySlice_l333_3 != 1'b0)) || (_zz_when_ArraySlice_l333_4 != 1'b0)) || (_zz_when_ArraySlice_l333_5 != 1'b0)) || (_zz_when_ArraySlice_l333_6 != 1'b0)) || (_zz_when_ArraySlice_l333_7 != 1'b0)));
  assign when_ArraySlice_l334 = (_zz_when_ArraySlice_l334 < _zz_when_ArraySlice_l334_1);
  assign _zz_19 = ({63'd0,1'b1} <<< selectWriteFifo);
  assign _zz_20 = ({63'd0,1'b1} <<< selectWriteFifo);
  assign _zz_io_push_valid_1 = inputStreamArrayData_valid;
  assign _zz_io_push_payload_1 = inputStreamArrayData_payload;
  assign inputStreamArrayData_fire_1 = (inputStreamArrayData_valid && inputStreamArrayData_ready);
  assign when_ArraySlice_l338 = ((_zz_when_ArraySlice_l338 == _zz_when_ArraySlice_l338_1) && inputStreamArrayData_fire_1);
  assign when_ArraySlice_l339 = (selectWriteFifo == _zz_when_ArraySlice_l339);
  always @(*) begin
    debug_0_50 = 1'b0;
    if(when_ArraySlice_l165_400) begin
      if(when_ArraySlice_l166_400) begin
        debug_0_50 = 1'b1;
      end else begin
        debug_0_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_400) begin
        debug_0_50 = 1'b1;
      end else begin
        debug_0_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_50 = 1'b0;
    if(when_ArraySlice_l165_401) begin
      if(when_ArraySlice_l166_401) begin
        debug_1_50 = 1'b1;
      end else begin
        debug_1_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_401) begin
        debug_1_50 = 1'b1;
      end else begin
        debug_1_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_50 = 1'b0;
    if(when_ArraySlice_l165_402) begin
      if(when_ArraySlice_l166_402) begin
        debug_2_50 = 1'b1;
      end else begin
        debug_2_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_402) begin
        debug_2_50 = 1'b1;
      end else begin
        debug_2_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_50 = 1'b0;
    if(when_ArraySlice_l165_403) begin
      if(when_ArraySlice_l166_403) begin
        debug_3_50 = 1'b1;
      end else begin
        debug_3_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_403) begin
        debug_3_50 = 1'b1;
      end else begin
        debug_3_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_50 = 1'b0;
    if(when_ArraySlice_l165_404) begin
      if(when_ArraySlice_l166_404) begin
        debug_4_50 = 1'b1;
      end else begin
        debug_4_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_404) begin
        debug_4_50 = 1'b1;
      end else begin
        debug_4_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_50 = 1'b0;
    if(when_ArraySlice_l165_405) begin
      if(when_ArraySlice_l166_405) begin
        debug_5_50 = 1'b1;
      end else begin
        debug_5_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_405) begin
        debug_5_50 = 1'b1;
      end else begin
        debug_5_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_50 = 1'b0;
    if(when_ArraySlice_l165_406) begin
      if(when_ArraySlice_l166_406) begin
        debug_6_50 = 1'b1;
      end else begin
        debug_6_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_406) begin
        debug_6_50 = 1'b1;
      end else begin
        debug_6_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_50 = 1'b0;
    if(when_ArraySlice_l165_407) begin
      if(when_ArraySlice_l166_407) begin
        debug_7_50 = 1'b1;
      end else begin
        debug_7_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_407) begin
        debug_7_50 = 1'b1;
      end else begin
        debug_7_50 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_400 = (_zz_when_ArraySlice_l165_400 <= selectWriteFifo);
  assign when_ArraySlice_l166_400 = (_zz_when_ArraySlice_l166_400 <= _zz_when_ArraySlice_l166_400_1);
  assign _zz_when_ArraySlice_l112_400 = (wReg % _zz__zz_when_ArraySlice_l112_400);
  assign when_ArraySlice_l112_400 = (_zz_when_ArraySlice_l112_400 != 6'h0);
  assign when_ArraySlice_l113_400 = (7'h40 <= _zz_when_ArraySlice_l113_400);
  always @(*) begin
    if(when_ArraySlice_l112_400) begin
      if(when_ArraySlice_l113_400) begin
        _zz_when_ArraySlice_l173_400 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_400 = (_zz__zz_when_ArraySlice_l173_400 - _zz__zz_when_ArraySlice_l173_400_3);
      end
    end else begin
      if(when_ArraySlice_l118_400) begin
        _zz_when_ArraySlice_l173_400 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_400 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_400 = (_zz_when_ArraySlice_l118_400 <= wReg);
  assign when_ArraySlice_l173_400 = (_zz_when_ArraySlice_l173_400_1 <= _zz_when_ArraySlice_l173_400_2);
  assign when_ArraySlice_l165_401 = (_zz_when_ArraySlice_l165_401 <= selectWriteFifo);
  assign when_ArraySlice_l166_401 = (_zz_when_ArraySlice_l166_401 <= _zz_when_ArraySlice_l166_401_1);
  assign _zz_when_ArraySlice_l112_401 = (wReg % _zz__zz_when_ArraySlice_l112_401);
  assign when_ArraySlice_l112_401 = (_zz_when_ArraySlice_l112_401 != 6'h0);
  assign when_ArraySlice_l113_401 = (7'h40 <= _zz_when_ArraySlice_l113_401);
  always @(*) begin
    if(when_ArraySlice_l112_401) begin
      if(when_ArraySlice_l113_401) begin
        _zz_when_ArraySlice_l173_401 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_401 = (_zz__zz_when_ArraySlice_l173_401 - _zz__zz_when_ArraySlice_l173_401_3);
      end
    end else begin
      if(when_ArraySlice_l118_401) begin
        _zz_when_ArraySlice_l173_401 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_401 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_401 = (_zz_when_ArraySlice_l118_401 <= wReg);
  assign when_ArraySlice_l173_401 = (_zz_when_ArraySlice_l173_401_1 <= _zz_when_ArraySlice_l173_401_3);
  assign when_ArraySlice_l165_402 = (_zz_when_ArraySlice_l165_402 <= selectWriteFifo);
  assign when_ArraySlice_l166_402 = (_zz_when_ArraySlice_l166_402 <= _zz_when_ArraySlice_l166_402_1);
  assign _zz_when_ArraySlice_l112_402 = (wReg % _zz__zz_when_ArraySlice_l112_402);
  assign when_ArraySlice_l112_402 = (_zz_when_ArraySlice_l112_402 != 6'h0);
  assign when_ArraySlice_l113_402 = (7'h40 <= _zz_when_ArraySlice_l113_402);
  always @(*) begin
    if(when_ArraySlice_l112_402) begin
      if(when_ArraySlice_l113_402) begin
        _zz_when_ArraySlice_l173_402 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_402 = (_zz__zz_when_ArraySlice_l173_402 - _zz__zz_when_ArraySlice_l173_402_3);
      end
    end else begin
      if(when_ArraySlice_l118_402) begin
        _zz_when_ArraySlice_l173_402 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_402 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_402 = (_zz_when_ArraySlice_l118_402 <= wReg);
  assign when_ArraySlice_l173_402 = (_zz_when_ArraySlice_l173_402_1 <= _zz_when_ArraySlice_l173_402_3);
  assign when_ArraySlice_l165_403 = (_zz_when_ArraySlice_l165_403 <= selectWriteFifo);
  assign when_ArraySlice_l166_403 = (_zz_when_ArraySlice_l166_403 <= _zz_when_ArraySlice_l166_403_1);
  assign _zz_when_ArraySlice_l112_403 = (wReg % _zz__zz_when_ArraySlice_l112_403);
  assign when_ArraySlice_l112_403 = (_zz_when_ArraySlice_l112_403 != 6'h0);
  assign when_ArraySlice_l113_403 = (7'h40 <= _zz_when_ArraySlice_l113_403);
  always @(*) begin
    if(when_ArraySlice_l112_403) begin
      if(when_ArraySlice_l113_403) begin
        _zz_when_ArraySlice_l173_403 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_403 = (_zz__zz_when_ArraySlice_l173_403 - _zz__zz_when_ArraySlice_l173_403_3);
      end
    end else begin
      if(when_ArraySlice_l118_403) begin
        _zz_when_ArraySlice_l173_403 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_403 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_403 = (_zz_when_ArraySlice_l118_403 <= wReg);
  assign when_ArraySlice_l173_403 = (_zz_when_ArraySlice_l173_403_1 <= _zz_when_ArraySlice_l173_403_3);
  assign when_ArraySlice_l165_404 = (_zz_when_ArraySlice_l165_404 <= selectWriteFifo);
  assign when_ArraySlice_l166_404 = (_zz_when_ArraySlice_l166_404 <= _zz_when_ArraySlice_l166_404_1);
  assign _zz_when_ArraySlice_l112_404 = (wReg % _zz__zz_when_ArraySlice_l112_404);
  assign when_ArraySlice_l112_404 = (_zz_when_ArraySlice_l112_404 != 6'h0);
  assign when_ArraySlice_l113_404 = (7'h40 <= _zz_when_ArraySlice_l113_404);
  always @(*) begin
    if(when_ArraySlice_l112_404) begin
      if(when_ArraySlice_l113_404) begin
        _zz_when_ArraySlice_l173_404 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_404 = (_zz__zz_when_ArraySlice_l173_404 - _zz__zz_when_ArraySlice_l173_404_3);
      end
    end else begin
      if(when_ArraySlice_l118_404) begin
        _zz_when_ArraySlice_l173_404 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_404 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_404 = (_zz_when_ArraySlice_l118_404 <= wReg);
  assign when_ArraySlice_l173_404 = (_zz_when_ArraySlice_l173_404_1 <= _zz_when_ArraySlice_l173_404_3);
  assign when_ArraySlice_l165_405 = (_zz_when_ArraySlice_l165_405 <= selectWriteFifo);
  assign when_ArraySlice_l166_405 = (_zz_when_ArraySlice_l166_405 <= _zz_when_ArraySlice_l166_405_2);
  assign _zz_when_ArraySlice_l112_405 = (wReg % _zz__zz_when_ArraySlice_l112_405);
  assign when_ArraySlice_l112_405 = (_zz_when_ArraySlice_l112_405 != 6'h0);
  assign when_ArraySlice_l113_405 = (7'h40 <= _zz_when_ArraySlice_l113_405);
  always @(*) begin
    if(when_ArraySlice_l112_405) begin
      if(when_ArraySlice_l113_405) begin
        _zz_when_ArraySlice_l173_405 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_405 = (_zz__zz_when_ArraySlice_l173_405 - _zz__zz_when_ArraySlice_l173_405_3);
      end
    end else begin
      if(when_ArraySlice_l118_405) begin
        _zz_when_ArraySlice_l173_405 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_405 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_405 = (_zz_when_ArraySlice_l118_405 <= wReg);
  assign when_ArraySlice_l173_405 = (_zz_when_ArraySlice_l173_405_1 <= _zz_when_ArraySlice_l173_405_3);
  assign when_ArraySlice_l165_406 = (_zz_when_ArraySlice_l165_406 <= selectWriteFifo);
  assign when_ArraySlice_l166_406 = (_zz_when_ArraySlice_l166_406 <= _zz_when_ArraySlice_l166_406_2);
  assign _zz_when_ArraySlice_l112_406 = (wReg % _zz__zz_when_ArraySlice_l112_406);
  assign when_ArraySlice_l112_406 = (_zz_when_ArraySlice_l112_406 != 6'h0);
  assign when_ArraySlice_l113_406 = (7'h40 <= _zz_when_ArraySlice_l113_406);
  always @(*) begin
    if(when_ArraySlice_l112_406) begin
      if(when_ArraySlice_l113_406) begin
        _zz_when_ArraySlice_l173_406 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_406 = (_zz__zz_when_ArraySlice_l173_406 - _zz__zz_when_ArraySlice_l173_406_3);
      end
    end else begin
      if(when_ArraySlice_l118_406) begin
        _zz_when_ArraySlice_l173_406 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_406 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_406 = (_zz_when_ArraySlice_l118_406 <= wReg);
  assign when_ArraySlice_l173_406 = (_zz_when_ArraySlice_l173_406_1 <= _zz_when_ArraySlice_l173_406_3);
  assign when_ArraySlice_l165_407 = (_zz_when_ArraySlice_l165_407 <= selectWriteFifo);
  assign when_ArraySlice_l166_407 = (_zz_when_ArraySlice_l166_407 <= _zz_when_ArraySlice_l166_407_2);
  assign _zz_when_ArraySlice_l112_407 = (wReg % _zz__zz_when_ArraySlice_l112_407);
  assign when_ArraySlice_l112_407 = (_zz_when_ArraySlice_l112_407 != 6'h0);
  assign when_ArraySlice_l113_407 = (7'h40 <= _zz_when_ArraySlice_l113_407);
  always @(*) begin
    if(when_ArraySlice_l112_407) begin
      if(when_ArraySlice_l113_407) begin
        _zz_when_ArraySlice_l173_407 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_407 = (_zz__zz_when_ArraySlice_l173_407 - _zz__zz_when_ArraySlice_l173_407_3);
      end
    end else begin
      if(when_ArraySlice_l118_407) begin
        _zz_when_ArraySlice_l173_407 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_407 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_407 = (_zz_when_ArraySlice_l118_407 <= wReg);
  assign when_ArraySlice_l173_407 = (_zz_when_ArraySlice_l173_407_1 <= _zz_when_ArraySlice_l173_407_3);
  assign when_ArraySlice_l350 = ((((((_zz_when_ArraySlice_l350 && _zz_when_ArraySlice_l350_1) && (holdReadOp_4 == _zz_when_ArraySlice_l350_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l350_3 && _zz_when_ArraySlice_l350_4) && (debug_4_50 == _zz_when_ArraySlice_l350_5)) && (debug_5_50 == 1'b1)) && (debug_6_50 == 1'b1)) && (debug_7_50 == 1'b1)));
  always @(*) begin
    debug_0_51 = 1'b0;
    if(when_ArraySlice_l165_408) begin
      if(when_ArraySlice_l166_408) begin
        debug_0_51 = 1'b1;
      end else begin
        debug_0_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_408) begin
        debug_0_51 = 1'b1;
      end else begin
        debug_0_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_51 = 1'b0;
    if(when_ArraySlice_l165_409) begin
      if(when_ArraySlice_l166_409) begin
        debug_1_51 = 1'b1;
      end else begin
        debug_1_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_409) begin
        debug_1_51 = 1'b1;
      end else begin
        debug_1_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_51 = 1'b0;
    if(when_ArraySlice_l165_410) begin
      if(when_ArraySlice_l166_410) begin
        debug_2_51 = 1'b1;
      end else begin
        debug_2_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_410) begin
        debug_2_51 = 1'b1;
      end else begin
        debug_2_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_51 = 1'b0;
    if(when_ArraySlice_l165_411) begin
      if(when_ArraySlice_l166_411) begin
        debug_3_51 = 1'b1;
      end else begin
        debug_3_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_411) begin
        debug_3_51 = 1'b1;
      end else begin
        debug_3_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_51 = 1'b0;
    if(when_ArraySlice_l165_412) begin
      if(when_ArraySlice_l166_412) begin
        debug_4_51 = 1'b1;
      end else begin
        debug_4_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_412) begin
        debug_4_51 = 1'b1;
      end else begin
        debug_4_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_51 = 1'b0;
    if(when_ArraySlice_l165_413) begin
      if(when_ArraySlice_l166_413) begin
        debug_5_51 = 1'b1;
      end else begin
        debug_5_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_413) begin
        debug_5_51 = 1'b1;
      end else begin
        debug_5_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_51 = 1'b0;
    if(when_ArraySlice_l165_414) begin
      if(when_ArraySlice_l166_414) begin
        debug_6_51 = 1'b1;
      end else begin
        debug_6_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_414) begin
        debug_6_51 = 1'b1;
      end else begin
        debug_6_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_51 = 1'b0;
    if(when_ArraySlice_l165_415) begin
      if(when_ArraySlice_l166_415) begin
        debug_7_51 = 1'b1;
      end else begin
        debug_7_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l173_415) begin
        debug_7_51 = 1'b1;
      end else begin
        debug_7_51 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l165_408 = (_zz_when_ArraySlice_l165_408 <= selectWriteFifo);
  assign when_ArraySlice_l166_408 = (_zz_when_ArraySlice_l166_408 <= _zz_when_ArraySlice_l166_408_1);
  assign _zz_when_ArraySlice_l112_408 = (wReg % _zz__zz_when_ArraySlice_l112_408);
  assign when_ArraySlice_l112_408 = (_zz_when_ArraySlice_l112_408 != 6'h0);
  assign when_ArraySlice_l113_408 = (7'h40 <= _zz_when_ArraySlice_l113_408);
  always @(*) begin
    if(when_ArraySlice_l112_408) begin
      if(when_ArraySlice_l113_408) begin
        _zz_when_ArraySlice_l173_408 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_408 = (_zz__zz_when_ArraySlice_l173_408 - _zz__zz_when_ArraySlice_l173_408_3);
      end
    end else begin
      if(when_ArraySlice_l118_408) begin
        _zz_when_ArraySlice_l173_408 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_408 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_408 = (_zz_when_ArraySlice_l118_408 <= wReg);
  assign when_ArraySlice_l173_408 = (_zz_when_ArraySlice_l173_408_1 <= _zz_when_ArraySlice_l173_408_2);
  assign when_ArraySlice_l165_409 = (_zz_when_ArraySlice_l165_409 <= selectWriteFifo);
  assign when_ArraySlice_l166_409 = (_zz_when_ArraySlice_l166_409 <= _zz_when_ArraySlice_l166_409_1);
  assign _zz_when_ArraySlice_l112_409 = (wReg % _zz__zz_when_ArraySlice_l112_409);
  assign when_ArraySlice_l112_409 = (_zz_when_ArraySlice_l112_409 != 6'h0);
  assign when_ArraySlice_l113_409 = (7'h40 <= _zz_when_ArraySlice_l113_409);
  always @(*) begin
    if(when_ArraySlice_l112_409) begin
      if(when_ArraySlice_l113_409) begin
        _zz_when_ArraySlice_l173_409 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_409 = (_zz__zz_when_ArraySlice_l173_409 - _zz__zz_when_ArraySlice_l173_409_3);
      end
    end else begin
      if(when_ArraySlice_l118_409) begin
        _zz_when_ArraySlice_l173_409 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_409 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_409 = (_zz_when_ArraySlice_l118_409 <= wReg);
  assign when_ArraySlice_l173_409 = (_zz_when_ArraySlice_l173_409_1 <= _zz_when_ArraySlice_l173_409_3);
  assign when_ArraySlice_l165_410 = (_zz_when_ArraySlice_l165_410 <= selectWriteFifo);
  assign when_ArraySlice_l166_410 = (_zz_when_ArraySlice_l166_410 <= _zz_when_ArraySlice_l166_410_1);
  assign _zz_when_ArraySlice_l112_410 = (wReg % _zz__zz_when_ArraySlice_l112_410);
  assign when_ArraySlice_l112_410 = (_zz_when_ArraySlice_l112_410 != 6'h0);
  assign when_ArraySlice_l113_410 = (7'h40 <= _zz_when_ArraySlice_l113_410);
  always @(*) begin
    if(when_ArraySlice_l112_410) begin
      if(when_ArraySlice_l113_410) begin
        _zz_when_ArraySlice_l173_410 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_410 = (_zz__zz_when_ArraySlice_l173_410 - _zz__zz_when_ArraySlice_l173_410_3);
      end
    end else begin
      if(when_ArraySlice_l118_410) begin
        _zz_when_ArraySlice_l173_410 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_410 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_410 = (_zz_when_ArraySlice_l118_410 <= wReg);
  assign when_ArraySlice_l173_410 = (_zz_when_ArraySlice_l173_410_1 <= _zz_when_ArraySlice_l173_410_3);
  assign when_ArraySlice_l165_411 = (_zz_when_ArraySlice_l165_411 <= selectWriteFifo);
  assign when_ArraySlice_l166_411 = (_zz_when_ArraySlice_l166_411 <= _zz_when_ArraySlice_l166_411_1);
  assign _zz_when_ArraySlice_l112_411 = (wReg % _zz__zz_when_ArraySlice_l112_411);
  assign when_ArraySlice_l112_411 = (_zz_when_ArraySlice_l112_411 != 6'h0);
  assign when_ArraySlice_l113_411 = (7'h40 <= _zz_when_ArraySlice_l113_411);
  always @(*) begin
    if(when_ArraySlice_l112_411) begin
      if(when_ArraySlice_l113_411) begin
        _zz_when_ArraySlice_l173_411 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_411 = (_zz__zz_when_ArraySlice_l173_411 - _zz__zz_when_ArraySlice_l173_411_3);
      end
    end else begin
      if(when_ArraySlice_l118_411) begin
        _zz_when_ArraySlice_l173_411 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_411 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_411 = (_zz_when_ArraySlice_l118_411 <= wReg);
  assign when_ArraySlice_l173_411 = (_zz_when_ArraySlice_l173_411_1 <= _zz_when_ArraySlice_l173_411_3);
  assign when_ArraySlice_l165_412 = (_zz_when_ArraySlice_l165_412 <= selectWriteFifo);
  assign when_ArraySlice_l166_412 = (_zz_when_ArraySlice_l166_412 <= _zz_when_ArraySlice_l166_412_1);
  assign _zz_when_ArraySlice_l112_412 = (wReg % _zz__zz_when_ArraySlice_l112_412);
  assign when_ArraySlice_l112_412 = (_zz_when_ArraySlice_l112_412 != 6'h0);
  assign when_ArraySlice_l113_412 = (7'h40 <= _zz_when_ArraySlice_l113_412);
  always @(*) begin
    if(when_ArraySlice_l112_412) begin
      if(when_ArraySlice_l113_412) begin
        _zz_when_ArraySlice_l173_412 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_412 = (_zz__zz_when_ArraySlice_l173_412 - _zz__zz_when_ArraySlice_l173_412_3);
      end
    end else begin
      if(when_ArraySlice_l118_412) begin
        _zz_when_ArraySlice_l173_412 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_412 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_412 = (_zz_when_ArraySlice_l118_412 <= wReg);
  assign when_ArraySlice_l173_412 = (_zz_when_ArraySlice_l173_412_1 <= _zz_when_ArraySlice_l173_412_3);
  assign when_ArraySlice_l165_413 = (_zz_when_ArraySlice_l165_413 <= selectWriteFifo);
  assign when_ArraySlice_l166_413 = (_zz_when_ArraySlice_l166_413 <= _zz_when_ArraySlice_l166_413_2);
  assign _zz_when_ArraySlice_l112_413 = (wReg % _zz__zz_when_ArraySlice_l112_413);
  assign when_ArraySlice_l112_413 = (_zz_when_ArraySlice_l112_413 != 6'h0);
  assign when_ArraySlice_l113_413 = (7'h40 <= _zz_when_ArraySlice_l113_413);
  always @(*) begin
    if(when_ArraySlice_l112_413) begin
      if(when_ArraySlice_l113_413) begin
        _zz_when_ArraySlice_l173_413 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_413 = (_zz__zz_when_ArraySlice_l173_413 - _zz__zz_when_ArraySlice_l173_413_3);
      end
    end else begin
      if(when_ArraySlice_l118_413) begin
        _zz_when_ArraySlice_l173_413 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_413 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_413 = (_zz_when_ArraySlice_l118_413 <= wReg);
  assign when_ArraySlice_l173_413 = (_zz_when_ArraySlice_l173_413_1 <= _zz_when_ArraySlice_l173_413_3);
  assign when_ArraySlice_l165_414 = (_zz_when_ArraySlice_l165_414 <= selectWriteFifo);
  assign when_ArraySlice_l166_414 = (_zz_when_ArraySlice_l166_414 <= _zz_when_ArraySlice_l166_414_2);
  assign _zz_when_ArraySlice_l112_414 = (wReg % _zz__zz_when_ArraySlice_l112_414);
  assign when_ArraySlice_l112_414 = (_zz_when_ArraySlice_l112_414 != 6'h0);
  assign when_ArraySlice_l113_414 = (7'h40 <= _zz_when_ArraySlice_l113_414);
  always @(*) begin
    if(when_ArraySlice_l112_414) begin
      if(when_ArraySlice_l113_414) begin
        _zz_when_ArraySlice_l173_414 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_414 = (_zz__zz_when_ArraySlice_l173_414 - _zz__zz_when_ArraySlice_l173_414_3);
      end
    end else begin
      if(when_ArraySlice_l118_414) begin
        _zz_when_ArraySlice_l173_414 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_414 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_414 = (_zz_when_ArraySlice_l118_414 <= wReg);
  assign when_ArraySlice_l173_414 = (_zz_when_ArraySlice_l173_414_1 <= _zz_when_ArraySlice_l173_414_3);
  assign when_ArraySlice_l165_415 = (_zz_when_ArraySlice_l165_415 <= selectWriteFifo);
  assign when_ArraySlice_l166_415 = (_zz_when_ArraySlice_l166_415 <= _zz_when_ArraySlice_l166_415_2);
  assign _zz_when_ArraySlice_l112_415 = (wReg % _zz__zz_when_ArraySlice_l112_415);
  assign when_ArraySlice_l112_415 = (_zz_when_ArraySlice_l112_415 != 6'h0);
  assign when_ArraySlice_l113_415 = (7'h40 <= _zz_when_ArraySlice_l113_415);
  always @(*) begin
    if(when_ArraySlice_l112_415) begin
      if(when_ArraySlice_l113_415) begin
        _zz_when_ArraySlice_l173_415 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_415 = (_zz__zz_when_ArraySlice_l173_415 - _zz__zz_when_ArraySlice_l173_415_3);
      end
    end else begin
      if(when_ArraySlice_l118_415) begin
        _zz_when_ArraySlice_l173_415 = 7'h40;
      end else begin
        _zz_when_ArraySlice_l173_415 = {1'd0, wReg};
      end
    end
  end

  assign when_ArraySlice_l118_415 = (_zz_when_ArraySlice_l118_415 <= wReg);
  assign when_ArraySlice_l173_415 = (_zz_when_ArraySlice_l173_415_1 <= _zz_when_ArraySlice_l173_415_3);
  assign when_ArraySlice_l189_8 = (selectWriteFifo == _zz_when_ArraySlice_l189_8);
  assign when_ArraySlice_l190_8 = (writeAround ^ readAround_0);
  always @(*) begin
    if(when_ArraySlice_l189_8) begin
      if(when_ArraySlice_l190_8) begin
        _zz_when_ArraySlice_l354 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l354 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l354 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_9 = (selectWriteFifo == _zz_when_ArraySlice_l189_9);
  assign when_ArraySlice_l190_9 = (writeAround ^ readAround_1);
  always @(*) begin
    if(when_ArraySlice_l189_9) begin
      if(when_ArraySlice_l190_9) begin
        _zz_when_ArraySlice_l354_1 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l354_1 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l354_1 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_10 = (selectWriteFifo == _zz_when_ArraySlice_l189_10);
  assign when_ArraySlice_l190_10 = (writeAround ^ readAround_2);
  always @(*) begin
    if(when_ArraySlice_l189_10) begin
      if(when_ArraySlice_l190_10) begin
        _zz_when_ArraySlice_l354_2 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l354_2 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l354_2 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_11 = (selectWriteFifo == _zz_when_ArraySlice_l189_11);
  assign when_ArraySlice_l190_11 = (writeAround ^ readAround_3);
  always @(*) begin
    if(when_ArraySlice_l189_11) begin
      if(when_ArraySlice_l190_11) begin
        _zz_when_ArraySlice_l354_3 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l354_3 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l354_3 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_12 = (selectWriteFifo == _zz_when_ArraySlice_l189_12);
  assign when_ArraySlice_l190_12 = (writeAround ^ readAround_4);
  always @(*) begin
    if(when_ArraySlice_l189_12) begin
      if(when_ArraySlice_l190_12) begin
        _zz_when_ArraySlice_l354_4 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l354_4 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l354_4 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_13 = (selectWriteFifo == _zz_when_ArraySlice_l189_13);
  assign when_ArraySlice_l190_13 = (writeAround ^ readAround_5);
  always @(*) begin
    if(when_ArraySlice_l189_13) begin
      if(when_ArraySlice_l190_13) begin
        _zz_when_ArraySlice_l354_5 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l354_5 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l354_5 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_14 = (selectWriteFifo == _zz_when_ArraySlice_l189_14);
  assign when_ArraySlice_l190_14 = (writeAround ^ readAround_6);
  always @(*) begin
    if(when_ArraySlice_l189_14) begin
      if(when_ArraySlice_l190_14) begin
        _zz_when_ArraySlice_l354_6 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l354_6 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l354_6 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_15 = (selectWriteFifo == _zz_when_ArraySlice_l189_15);
  assign when_ArraySlice_l190_15 = (writeAround ^ readAround_7);
  always @(*) begin
    if(when_ArraySlice_l189_15) begin
      if(when_ArraySlice_l190_15) begin
        _zz_when_ArraySlice_l354_7 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l354_7 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l354_7 = 1'b0;
    end
  end

  assign when_ArraySlice_l354 = (((((_zz_when_ArraySlice_l354_8 && _zz_when_ArraySlice_l354_12) && (holdReadOp_6 == _zz_when_ArraySlice_l354_13)) && (holdReadOp_7 == 1'b1)) && (! ((_zz_when_ArraySlice_l354_14 && _zz_when_ArraySlice_l354_18) && (debug_7_51 == _zz_when_ArraySlice_l354_19)))) && (! (((_zz_when_ArraySlice_l354_20 || _zz_when_ArraySlice_l354_24) || (_zz_when_ArraySlice_l354_6 != _zz_when_ArraySlice_l354_25)) || (_zz_when_ArraySlice_l354_7 != 1'b0))));
  assign when_ArraySlice_l189_16 = (selectWriteFifo == _zz_when_ArraySlice_l189_16);
  assign when_ArraySlice_l190_16 = (writeAround ^ readAround_0);
  always @(*) begin
    if(when_ArraySlice_l189_16) begin
      if(when_ArraySlice_l190_16) begin
        _zz_when_ArraySlice_l358 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l358 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l358 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_17 = (selectWriteFifo == _zz_when_ArraySlice_l189_17);
  assign when_ArraySlice_l190_17 = (writeAround ^ readAround_1);
  always @(*) begin
    if(when_ArraySlice_l189_17) begin
      if(when_ArraySlice_l190_17) begin
        _zz_when_ArraySlice_l358_1 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l358_1 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l358_1 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_18 = (selectWriteFifo == _zz_when_ArraySlice_l189_18);
  assign when_ArraySlice_l190_18 = (writeAround ^ readAround_2);
  always @(*) begin
    if(when_ArraySlice_l189_18) begin
      if(when_ArraySlice_l190_18) begin
        _zz_when_ArraySlice_l358_2 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l358_2 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l358_2 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_19 = (selectWriteFifo == _zz_when_ArraySlice_l189_19);
  assign when_ArraySlice_l190_19 = (writeAround ^ readAround_3);
  always @(*) begin
    if(when_ArraySlice_l189_19) begin
      if(when_ArraySlice_l190_19) begin
        _zz_when_ArraySlice_l358_3 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l358_3 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l358_3 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_20 = (selectWriteFifo == _zz_when_ArraySlice_l189_20);
  assign when_ArraySlice_l190_20 = (writeAround ^ readAround_4);
  always @(*) begin
    if(when_ArraySlice_l189_20) begin
      if(when_ArraySlice_l190_20) begin
        _zz_when_ArraySlice_l358_4 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l358_4 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l358_4 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_21 = (selectWriteFifo == _zz_when_ArraySlice_l189_21);
  assign when_ArraySlice_l190_21 = (writeAround ^ readAround_5);
  always @(*) begin
    if(when_ArraySlice_l189_21) begin
      if(when_ArraySlice_l190_21) begin
        _zz_when_ArraySlice_l358_5 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l358_5 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l358_5 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_22 = (selectWriteFifo == _zz_when_ArraySlice_l189_22);
  assign when_ArraySlice_l190_22 = (writeAround ^ readAround_6);
  always @(*) begin
    if(when_ArraySlice_l189_22) begin
      if(when_ArraySlice_l190_22) begin
        _zz_when_ArraySlice_l358_6 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l358_6 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l358_6 = 1'b0;
    end
  end

  assign when_ArraySlice_l189_23 = (selectWriteFifo == _zz_when_ArraySlice_l189_23);
  assign when_ArraySlice_l190_23 = (writeAround ^ readAround_7);
  always @(*) begin
    if(when_ArraySlice_l189_23) begin
      if(when_ArraySlice_l190_23) begin
        _zz_when_ArraySlice_l358_7 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l358_7 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l358_7 = 1'b0;
    end
  end

  assign when_ArraySlice_l358 = ((((((((_zz_when_ArraySlice_l358 != 1'b0) || (_zz_when_ArraySlice_l358_1 != 1'b0)) || (_zz_when_ArraySlice_l358_2 != 1'b0)) || (_zz_when_ArraySlice_l358_3 != 1'b0)) || (_zz_when_ArraySlice_l358_4 != 1'b0)) || (_zz_when_ArraySlice_l358_5 != 1'b0)) || (_zz_when_ArraySlice_l358_6 != 1'b0)) || (_zz_when_ArraySlice_l358_7 != 1'b0));
  assign when_ArraySlice_l361 = (! allowPadding_0);
  assign when_ArraySlice_l361_1 = (! allowPadding_1);
  assign when_ArraySlice_l361_2 = (! allowPadding_2);
  assign when_ArraySlice_l361_3 = (! allowPadding_3);
  assign when_ArraySlice_l361_4 = (! allowPadding_4);
  assign when_ArraySlice_l361_5 = (! allowPadding_5);
  assign when_ArraySlice_l361_6 = (! allowPadding_6);
  assign when_ArraySlice_l361_7 = (! allowPadding_7);
  assign stateIndicate = arraySliceStateMachine_stateReg;
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      wReg <= 6'h3f;
      hReg <= 6'h3f;
      aReg <= 3'b111;
      bReg <= 3'b111;
      handshakeTimes_0_value <= 13'h0;
      handshakeTimes_1_value <= 13'h0;
      handshakeTimes_2_value <= 13'h0;
      handshakeTimes_3_value <= 13'h0;
      handshakeTimes_4_value <= 13'h0;
      handshakeTimes_5_value <= 13'h0;
      handshakeTimes_6_value <= 13'h0;
      handshakeTimes_7_value <= 13'h0;
      selectWriteFifo <= 6'h0;
      selectReadFifo_0 <= 6'h0;
      selectReadFifo_1 <= 6'h0;
      selectReadFifo_2 <= 6'h0;
      selectReadFifo_3 <= 6'h0;
      selectReadFifo_4 <= 6'h0;
      selectReadFifo_5 <= 6'h0;
      selectReadFifo_6 <= 6'h0;
      selectReadFifo_7 <= 6'h0;
      holdReadOp_0 <= 1'b0;
      holdReadOp_1 <= 1'b0;
      holdReadOp_2 <= 1'b0;
      holdReadOp_3 <= 1'b0;
      holdReadOp_4 <= 1'b0;
      holdReadOp_5 <= 1'b0;
      holdReadOp_6 <= 1'b0;
      holdReadOp_7 <= 1'b0;
      allowPadding_0 <= 1'b1;
      allowPadding_1 <= 1'b1;
      allowPadding_2 <= 1'b1;
      allowPadding_3 <= 1'b1;
      allowPadding_4 <= 1'b1;
      allowPadding_5 <= 1'b1;
      allowPadding_6 <= 1'b1;
      allowPadding_7 <= 1'b1;
      outSliceNumb_0_value <= 7'h0;
      outSliceNumb_1_value <= 7'h0;
      outSliceNumb_2_value <= 7'h0;
      outSliceNumb_3_value <= 7'h0;
      outSliceNumb_4_value <= 7'h0;
      outSliceNumb_5_value <= 7'h0;
      outSliceNumb_6_value <= 7'h0;
      outSliceNumb_7_value <= 7'h0;
      writeAround <= 1'b0;
      readAround_0 <= 1'b0;
      readAround_1 <= 1'b0;
      readAround_2 <= 1'b0;
      readAround_3 <= 1'b0;
      readAround_4 <= 1'b0;
      readAround_5 <= 1'b0;
      readAround_6 <= 1'b0;
      readAround_7 <= 1'b0;
      arraySliceStateMachine_stateReg <= arraySliceStateMachine_enumDef_BOOT;
    end else begin
      wReg <= inputFeatureMapWidth;
      hReg <= inputFeatureMapHeight;
      aReg <= outputFeatureMapHeight;
      bReg <= outputFeatureMapWidth;
      handshakeTimes_0_value <= handshakeTimes_0_valueNext;
      handshakeTimes_1_value <= handshakeTimes_1_valueNext;
      handshakeTimes_2_value <= handshakeTimes_2_valueNext;
      handshakeTimes_3_value <= handshakeTimes_3_valueNext;
      handshakeTimes_4_value <= handshakeTimes_4_valueNext;
      handshakeTimes_5_value <= handshakeTimes_5_valueNext;
      handshakeTimes_6_value <= handshakeTimes_6_valueNext;
      handshakeTimes_7_value <= handshakeTimes_7_valueNext;
      outSliceNumb_0_value <= outSliceNumb_0_valueNext;
      outSliceNumb_1_value <= outSliceNumb_1_valueNext;
      outSliceNumb_2_value <= outSliceNumb_2_valueNext;
      outSliceNumb_3_value <= outSliceNumb_3_valueNext;
      outSliceNumb_4_value <= outSliceNumb_4_valueNext;
      outSliceNumb_5_value <= outSliceNumb_5_valueNext;
      outSliceNumb_6_value <= outSliceNumb_6_valueNext;
      outSliceNumb_7_value <= outSliceNumb_7_valueNext;
      arraySliceStateMachine_stateReg <= arraySliceStateMachine_stateNext;
      case(arraySliceStateMachine_stateReg)
        arraySliceStateMachine_enumDef_writeDataOnly : begin
          if(when_ArraySlice_l215) begin
            if(when_ArraySlice_l216) begin
              selectWriteFifo <= 6'h0;
              writeAround <= (! writeAround);
            end else begin
              selectWriteFifo <= (selectWriteFifo + _zz_selectWriteFifo);
            end
          end
          if(when_ArraySlice_l223) begin
            if(holdReadOp_0) begin
              holdReadOp_0 <= 1'b0;
            end
            if(when_ArraySlice_l229) begin
              allowPadding_0 <= 1'b1;
            end
            if(holdReadOp_1) begin
              holdReadOp_1 <= 1'b0;
            end
            if(when_ArraySlice_l229_1) begin
              allowPadding_1 <= 1'b1;
            end
            if(holdReadOp_2) begin
              holdReadOp_2 <= 1'b0;
            end
            if(when_ArraySlice_l229_2) begin
              allowPadding_2 <= 1'b1;
            end
            if(holdReadOp_3) begin
              holdReadOp_3 <= 1'b0;
            end
            if(when_ArraySlice_l229_3) begin
              allowPadding_3 <= 1'b1;
            end
            if(holdReadOp_4) begin
              holdReadOp_4 <= 1'b0;
            end
            if(when_ArraySlice_l229_4) begin
              allowPadding_4 <= 1'b1;
            end
            if(holdReadOp_5) begin
              holdReadOp_5 <= 1'b0;
            end
            if(when_ArraySlice_l229_5) begin
              allowPadding_5 <= 1'b1;
            end
            if(holdReadOp_6) begin
              holdReadOp_6 <= 1'b0;
            end
            if(when_ArraySlice_l229_6) begin
              allowPadding_6 <= 1'b1;
            end
            if(holdReadOp_7) begin
              holdReadOp_7 <= 1'b0;
            end
            if(when_ArraySlice_l229_7) begin
              allowPadding_7 <= 1'b1;
            end
          end
        end
        arraySliceStateMachine_enumDef_readDataOnly : begin
          if(when_ArraySlice_l373) begin
            if(when_ArraySlice_l379) begin
              if(when_ArraySlice_l380) begin
                if(when_ArraySlice_l381) begin
                  selectReadFifo_0 <= (_zz_selectReadFifo_0 + _zz_selectReadFifo_0_2);
                end else begin
                  if(when_ArraySlice_l384) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + _zz_selectReadFifo_0_4);
                  end
                end
              end
              if(when_ArraySlice_l389) begin
                if(when_ArraySlice_l390) begin
                  if(when_ArraySlice_l392) begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_6 + _zz_selectReadFifo_0_8);
                  end else begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_10 + _zz_selectReadFifo_0_12);
                    if(when_ArraySlice_l398) begin
                      holdReadOp_0 <= 1'b1;
                    end
                    if(when_ArraySlice_l401) begin
                      allowPadding_0 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l405) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + _zz_selectReadFifo_0_14);
                  end
                end
              end
              if(when_ArraySlice_l409) begin
                if(when_ArraySlice_l410) begin
                  if(when_ArraySlice_l412) begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_16 + _zz_selectReadFifo_0_18);
                  end else begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_20 + _zz_selectReadFifo_0_22);
                    if(when_ArraySlice_l418) begin
                      holdReadOp_0 <= 1'b1;
                    end
                    if(when_ArraySlice_l421) begin
                      allowPadding_0 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l425) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + _zz_selectReadFifo_0_24);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l434) begin
              if(when_ArraySlice_l436) begin
                if(when_ArraySlice_l437) begin
                  selectReadFifo_0 <= (_zz_selectReadFifo_0_26 + _zz_selectReadFifo_0_28);
                end else begin
                  selectReadFifo_0 <= 6'h0;
                  readAround_0 <= (! readAround_0);
                  if(when_ArraySlice_l444) begin
                    holdReadOp_0 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l448) begin
                  selectReadFifo_0 <= (selectReadFifo_0 + _zz_selectReadFifo_0_30);
                end
              end
            end
          end
          if(when_ArraySlice_l373_1) begin
            if(when_ArraySlice_l379_1) begin
              if(when_ArraySlice_l380_1) begin
                if(when_ArraySlice_l381_1) begin
                  selectReadFifo_1 <= (_zz_selectReadFifo_1 + _zz_selectReadFifo_1_2);
                end else begin
                  if(when_ArraySlice_l384_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + _zz_selectReadFifo_1_4);
                  end
                end
              end
              if(when_ArraySlice_l389_1) begin
                if(when_ArraySlice_l390_1) begin
                  if(when_ArraySlice_l392_1) begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_6 + _zz_selectReadFifo_1_8);
                  end else begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_10 + _zz_selectReadFifo_1_12);
                    if(when_ArraySlice_l398_1) begin
                      holdReadOp_1 <= 1'b1;
                    end
                    if(when_ArraySlice_l401_1) begin
                      allowPadding_1 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l405_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + _zz_selectReadFifo_1_14);
                  end
                end
              end
              if(when_ArraySlice_l409_1) begin
                if(when_ArraySlice_l410_1) begin
                  if(when_ArraySlice_l412_1) begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_16 + _zz_selectReadFifo_1_18);
                  end else begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_20 + _zz_selectReadFifo_1_22);
                    if(when_ArraySlice_l418_1) begin
                      holdReadOp_1 <= 1'b1;
                    end
                    if(when_ArraySlice_l421_1) begin
                      allowPadding_1 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l425_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + _zz_selectReadFifo_1_24);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l434_1) begin
              if(when_ArraySlice_l436_1) begin
                if(when_ArraySlice_l437_1) begin
                  selectReadFifo_1 <= (_zz_selectReadFifo_1_26 + _zz_selectReadFifo_1_28);
                end else begin
                  selectReadFifo_1 <= 6'h0;
                  readAround_1 <= (! readAround_1);
                  if(when_ArraySlice_l444_1) begin
                    holdReadOp_1 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l448_1) begin
                  selectReadFifo_1 <= (selectReadFifo_1 + _zz_selectReadFifo_1_30);
                end
              end
            end
          end
          if(when_ArraySlice_l373_2) begin
            if(when_ArraySlice_l379_2) begin
              if(when_ArraySlice_l380_2) begin
                if(when_ArraySlice_l381_2) begin
                  selectReadFifo_2 <= (_zz_selectReadFifo_2 + _zz_selectReadFifo_2_2);
                end else begin
                  if(when_ArraySlice_l384_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + _zz_selectReadFifo_2_4);
                  end
                end
              end
              if(when_ArraySlice_l389_2) begin
                if(when_ArraySlice_l390_2) begin
                  if(when_ArraySlice_l392_2) begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_6 + _zz_selectReadFifo_2_8);
                  end else begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_10 + _zz_selectReadFifo_2_12);
                    if(when_ArraySlice_l398_2) begin
                      holdReadOp_2 <= 1'b1;
                    end
                    if(when_ArraySlice_l401_2) begin
                      allowPadding_2 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l405_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + _zz_selectReadFifo_2_14);
                  end
                end
              end
              if(when_ArraySlice_l409_2) begin
                if(when_ArraySlice_l410_2) begin
                  if(when_ArraySlice_l412_2) begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_16 + _zz_selectReadFifo_2_18);
                  end else begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_20 + _zz_selectReadFifo_2_22);
                    if(when_ArraySlice_l418_2) begin
                      holdReadOp_2 <= 1'b1;
                    end
                    if(when_ArraySlice_l421_2) begin
                      allowPadding_2 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l425_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + _zz_selectReadFifo_2_24);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l434_2) begin
              if(when_ArraySlice_l436_2) begin
                if(when_ArraySlice_l437_2) begin
                  selectReadFifo_2 <= (_zz_selectReadFifo_2_26 + _zz_selectReadFifo_2_28);
                end else begin
                  selectReadFifo_2 <= 6'h0;
                  readAround_2 <= (! readAround_2);
                  if(when_ArraySlice_l444_2) begin
                    holdReadOp_2 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l448_2) begin
                  selectReadFifo_2 <= (selectReadFifo_2 + _zz_selectReadFifo_2_30);
                end
              end
            end
          end
          if(when_ArraySlice_l373_3) begin
            if(when_ArraySlice_l379_3) begin
              if(when_ArraySlice_l380_3) begin
                if(when_ArraySlice_l381_3) begin
                  selectReadFifo_3 <= (_zz_selectReadFifo_3 + _zz_selectReadFifo_3_2);
                end else begin
                  if(when_ArraySlice_l384_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + _zz_selectReadFifo_3_4);
                  end
                end
              end
              if(when_ArraySlice_l389_3) begin
                if(when_ArraySlice_l390_3) begin
                  if(when_ArraySlice_l392_3) begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_6 + _zz_selectReadFifo_3_8);
                  end else begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_10 + _zz_selectReadFifo_3_12);
                    if(when_ArraySlice_l398_3) begin
                      holdReadOp_3 <= 1'b1;
                    end
                    if(when_ArraySlice_l401_3) begin
                      allowPadding_3 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l405_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + _zz_selectReadFifo_3_14);
                  end
                end
              end
              if(when_ArraySlice_l409_3) begin
                if(when_ArraySlice_l410_3) begin
                  if(when_ArraySlice_l412_3) begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_16 + _zz_selectReadFifo_3_18);
                  end else begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_20 + _zz_selectReadFifo_3_22);
                    if(when_ArraySlice_l418_3) begin
                      holdReadOp_3 <= 1'b1;
                    end
                    if(when_ArraySlice_l421_3) begin
                      allowPadding_3 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l425_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + _zz_selectReadFifo_3_24);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l434_3) begin
              if(when_ArraySlice_l436_3) begin
                if(when_ArraySlice_l437_3) begin
                  selectReadFifo_3 <= (_zz_selectReadFifo_3_26 + _zz_selectReadFifo_3_28);
                end else begin
                  selectReadFifo_3 <= 6'h0;
                  readAround_3 <= (! readAround_3);
                  if(when_ArraySlice_l444_3) begin
                    holdReadOp_3 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l448_3) begin
                  selectReadFifo_3 <= (selectReadFifo_3 + _zz_selectReadFifo_3_30);
                end
              end
            end
          end
          if(when_ArraySlice_l373_4) begin
            if(when_ArraySlice_l379_4) begin
              if(when_ArraySlice_l380_4) begin
                if(when_ArraySlice_l381_4) begin
                  selectReadFifo_4 <= (_zz_selectReadFifo_4 + _zz_selectReadFifo_4_2);
                end else begin
                  if(when_ArraySlice_l384_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + _zz_selectReadFifo_4_4);
                  end
                end
              end
              if(when_ArraySlice_l389_4) begin
                if(when_ArraySlice_l390_4) begin
                  if(when_ArraySlice_l392_4) begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_6 + _zz_selectReadFifo_4_8);
                  end else begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_10 + _zz_selectReadFifo_4_12);
                    if(when_ArraySlice_l398_4) begin
                      holdReadOp_4 <= 1'b1;
                    end
                    if(when_ArraySlice_l401_4) begin
                      allowPadding_4 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l405_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + _zz_selectReadFifo_4_14);
                  end
                end
              end
              if(when_ArraySlice_l409_4) begin
                if(when_ArraySlice_l410_4) begin
                  if(when_ArraySlice_l412_4) begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_16 + _zz_selectReadFifo_4_18);
                  end else begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_20 + _zz_selectReadFifo_4_22);
                    if(when_ArraySlice_l418_4) begin
                      holdReadOp_4 <= 1'b1;
                    end
                    if(when_ArraySlice_l421_4) begin
                      allowPadding_4 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l425_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + _zz_selectReadFifo_4_24);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l434_4) begin
              if(when_ArraySlice_l436_4) begin
                if(when_ArraySlice_l437_4) begin
                  selectReadFifo_4 <= (_zz_selectReadFifo_4_26 + _zz_selectReadFifo_4_28);
                end else begin
                  selectReadFifo_4 <= 6'h0;
                  readAround_4 <= (! readAround_4);
                  if(when_ArraySlice_l444_4) begin
                    holdReadOp_4 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l448_4) begin
                  selectReadFifo_4 <= (selectReadFifo_4 + _zz_selectReadFifo_4_30);
                end
              end
            end
          end
          if(when_ArraySlice_l373_5) begin
            if(when_ArraySlice_l379_5) begin
              if(when_ArraySlice_l380_5) begin
                if(when_ArraySlice_l381_5) begin
                  selectReadFifo_5 <= (_zz_selectReadFifo_5 + _zz_selectReadFifo_5_2);
                end else begin
                  if(when_ArraySlice_l384_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + _zz_selectReadFifo_5_4);
                  end
                end
              end
              if(when_ArraySlice_l389_5) begin
                if(when_ArraySlice_l390_5) begin
                  if(when_ArraySlice_l392_5) begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_6 + _zz_selectReadFifo_5_8);
                  end else begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_10 + _zz_selectReadFifo_5_12);
                    if(when_ArraySlice_l398_5) begin
                      holdReadOp_5 <= 1'b1;
                    end
                    if(when_ArraySlice_l401_5) begin
                      allowPadding_5 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l405_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + _zz_selectReadFifo_5_14);
                  end
                end
              end
              if(when_ArraySlice_l409_5) begin
                if(when_ArraySlice_l410_5) begin
                  if(when_ArraySlice_l412_5) begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_16 + _zz_selectReadFifo_5_18);
                  end else begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_20 + _zz_selectReadFifo_5_22);
                    if(when_ArraySlice_l418_5) begin
                      holdReadOp_5 <= 1'b1;
                    end
                    if(when_ArraySlice_l421_5) begin
                      allowPadding_5 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l425_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + _zz_selectReadFifo_5_24);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l434_5) begin
              if(when_ArraySlice_l436_5) begin
                if(when_ArraySlice_l437_5) begin
                  selectReadFifo_5 <= (_zz_selectReadFifo_5_26 + _zz_selectReadFifo_5_28);
                end else begin
                  selectReadFifo_5 <= 6'h0;
                  readAround_5 <= (! readAround_5);
                  if(when_ArraySlice_l444_5) begin
                    holdReadOp_5 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l448_5) begin
                  selectReadFifo_5 <= (selectReadFifo_5 + _zz_selectReadFifo_5_30);
                end
              end
            end
          end
          if(when_ArraySlice_l373_6) begin
            if(when_ArraySlice_l379_6) begin
              if(when_ArraySlice_l380_6) begin
                if(when_ArraySlice_l381_6) begin
                  selectReadFifo_6 <= (_zz_selectReadFifo_6 + _zz_selectReadFifo_6_2);
                end else begin
                  if(when_ArraySlice_l384_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + _zz_selectReadFifo_6_4);
                  end
                end
              end
              if(when_ArraySlice_l389_6) begin
                if(when_ArraySlice_l390_6) begin
                  if(when_ArraySlice_l392_6) begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_6 + _zz_selectReadFifo_6_8);
                  end else begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_10 + _zz_selectReadFifo_6_12);
                    if(when_ArraySlice_l398_6) begin
                      holdReadOp_6 <= 1'b1;
                    end
                    if(when_ArraySlice_l401_6) begin
                      allowPadding_6 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l405_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + _zz_selectReadFifo_6_14);
                  end
                end
              end
              if(when_ArraySlice_l409_6) begin
                if(when_ArraySlice_l410_6) begin
                  if(when_ArraySlice_l412_6) begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_16 + _zz_selectReadFifo_6_18);
                  end else begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_20 + _zz_selectReadFifo_6_22);
                    if(when_ArraySlice_l418_6) begin
                      holdReadOp_6 <= 1'b1;
                    end
                    if(when_ArraySlice_l421_6) begin
                      allowPadding_6 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l425_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + _zz_selectReadFifo_6_24);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l434_6) begin
              if(when_ArraySlice_l436_6) begin
                if(when_ArraySlice_l437_6) begin
                  selectReadFifo_6 <= (_zz_selectReadFifo_6_26 + _zz_selectReadFifo_6_28);
                end else begin
                  selectReadFifo_6 <= 6'h0;
                  readAround_6 <= (! readAround_6);
                  if(when_ArraySlice_l444_6) begin
                    holdReadOp_6 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l448_6) begin
                  selectReadFifo_6 <= (selectReadFifo_6 + _zz_selectReadFifo_6_30);
                end
              end
            end
          end
          if(when_ArraySlice_l373_7) begin
            if(when_ArraySlice_l379_7) begin
              if(when_ArraySlice_l380_7) begin
                if(when_ArraySlice_l381_7) begin
                  selectReadFifo_7 <= (_zz_selectReadFifo_7 + _zz_selectReadFifo_7_2);
                end else begin
                  if(when_ArraySlice_l384_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + _zz_selectReadFifo_7_4);
                  end
                end
              end
              if(when_ArraySlice_l389_7) begin
                if(when_ArraySlice_l390_7) begin
                  if(when_ArraySlice_l392_7) begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_6 + _zz_selectReadFifo_7_8);
                  end else begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_10 + _zz_selectReadFifo_7_12);
                    if(when_ArraySlice_l398_7) begin
                      holdReadOp_7 <= 1'b1;
                    end
                    if(when_ArraySlice_l401_7) begin
                      allowPadding_7 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l405_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + _zz_selectReadFifo_7_14);
                  end
                end
              end
              if(when_ArraySlice_l409_7) begin
                if(when_ArraySlice_l410_7) begin
                  if(when_ArraySlice_l412_7) begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_16 + _zz_selectReadFifo_7_18);
                  end else begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_20 + _zz_selectReadFifo_7_22);
                    if(when_ArraySlice_l418_7) begin
                      holdReadOp_7 <= 1'b1;
                    end
                    if(when_ArraySlice_l421_7) begin
                      allowPadding_7 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l425_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + _zz_selectReadFifo_7_24);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l434_7) begin
              if(when_ArraySlice_l436_7) begin
                if(when_ArraySlice_l437_7) begin
                  selectReadFifo_7 <= (_zz_selectReadFifo_7_26 + _zz_selectReadFifo_7_28);
                end else begin
                  selectReadFifo_7 <= 6'h0;
                  readAround_7 <= (! readAround_7);
                  if(when_ArraySlice_l444_7) begin
                    holdReadOp_7 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l448_7) begin
                  selectReadFifo_7 <= (selectReadFifo_7 + _zz_selectReadFifo_7_30);
                end
              end
            end
          end
          if(when_ArraySlice_l465) begin
            holdReadOp_0 <= 1'b0;
            if(when_ArraySlice_l468) begin
              allowPadding_0 <= 1'b1;
            end
            holdReadOp_1 <= 1'b0;
            if(when_ArraySlice_l468_1) begin
              allowPadding_1 <= 1'b1;
            end
            holdReadOp_2 <= 1'b0;
            if(when_ArraySlice_l468_2) begin
              allowPadding_2 <= 1'b1;
            end
            holdReadOp_3 <= 1'b0;
            if(when_ArraySlice_l468_3) begin
              allowPadding_3 <= 1'b1;
            end
            holdReadOp_4 <= 1'b0;
            if(when_ArraySlice_l468_4) begin
              allowPadding_4 <= 1'b1;
            end
            holdReadOp_5 <= 1'b0;
            if(when_ArraySlice_l468_5) begin
              allowPadding_5 <= 1'b1;
            end
            holdReadOp_6 <= 1'b0;
            if(when_ArraySlice_l468_6) begin
              allowPadding_6 <= 1'b1;
            end
            holdReadOp_7 <= 1'b0;
            if(when_ArraySlice_l468_7) begin
              allowPadding_7 <= 1'b1;
            end
          end
        end
        arraySliceStateMachine_enumDef_readWriteData : begin
          if(when_ArraySlice_l240) begin
            if(when_ArraySlice_l246) begin
              if(when_ArraySlice_l247) begin
                if(when_ArraySlice_l248) begin
                  selectReadFifo_0 <= (_zz_selectReadFifo_0_32 + _zz_selectReadFifo_0_34);
                end else begin
                  if(when_ArraySlice_l251) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + _zz_selectReadFifo_0_36);
                  end
                end
              end
              if(when_ArraySlice_l256) begin
                if(when_ArraySlice_l257) begin
                  if(when_ArraySlice_l259) begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_38 + _zz_selectReadFifo_0_40);
                  end else begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_42 + _zz_selectReadFifo_0_44);
                    if(when_ArraySlice_l265) begin
                      holdReadOp_0 <= 1'b1;
                    end
                    if(when_ArraySlice_l268) begin
                      allowPadding_0 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l272) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + _zz_selectReadFifo_0_46);
                  end
                end
              end
              if(when_ArraySlice_l276) begin
                if(when_ArraySlice_l277) begin
                  if(when_ArraySlice_l279) begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_48 + _zz_selectReadFifo_0_50);
                  end else begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_52 + _zz_selectReadFifo_0_54);
                    if(when_ArraySlice_l285) begin
                      holdReadOp_0 <= 1'b1;
                    end
                    if(when_ArraySlice_l288) begin
                      allowPadding_0 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l292) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + _zz_selectReadFifo_0_56);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l301) begin
              if(when_ArraySlice_l303) begin
                if(when_ArraySlice_l304) begin
                  selectReadFifo_0 <= (_zz_selectReadFifo_0_58 + _zz_selectReadFifo_0_60);
                end else begin
                  selectReadFifo_0 <= 6'h0;
                  readAround_0 <= (! readAround_0);
                  if(when_ArraySlice_l311) begin
                    holdReadOp_0 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l315) begin
                  selectReadFifo_0 <= (selectReadFifo_0 + _zz_selectReadFifo_0_62);
                end
              end
            end
          end
          if(when_ArraySlice_l240_1) begin
            if(when_ArraySlice_l246_1) begin
              if(when_ArraySlice_l247_1) begin
                if(when_ArraySlice_l248_1) begin
                  selectReadFifo_1 <= (_zz_selectReadFifo_1_32 + _zz_selectReadFifo_1_34);
                end else begin
                  if(when_ArraySlice_l251_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + _zz_selectReadFifo_1_36);
                  end
                end
              end
              if(when_ArraySlice_l256_1) begin
                if(when_ArraySlice_l257_1) begin
                  if(when_ArraySlice_l259_1) begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_38 + _zz_selectReadFifo_1_40);
                  end else begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_42 + _zz_selectReadFifo_1_44);
                    if(when_ArraySlice_l265_1) begin
                      holdReadOp_1 <= 1'b1;
                    end
                    if(when_ArraySlice_l268_1) begin
                      allowPadding_1 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l272_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + _zz_selectReadFifo_1_46);
                  end
                end
              end
              if(when_ArraySlice_l276_1) begin
                if(when_ArraySlice_l277_1) begin
                  if(when_ArraySlice_l279_1) begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_48 + _zz_selectReadFifo_1_50);
                  end else begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_52 + _zz_selectReadFifo_1_54);
                    if(when_ArraySlice_l285_1) begin
                      holdReadOp_1 <= 1'b1;
                    end
                    if(when_ArraySlice_l288_1) begin
                      allowPadding_1 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l292_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + _zz_selectReadFifo_1_56);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l301_1) begin
              if(when_ArraySlice_l303_1) begin
                if(when_ArraySlice_l304_1) begin
                  selectReadFifo_1 <= (_zz_selectReadFifo_1_58 + _zz_selectReadFifo_1_60);
                end else begin
                  selectReadFifo_1 <= 6'h0;
                  readAround_1 <= (! readAround_1);
                  if(when_ArraySlice_l311_1) begin
                    holdReadOp_1 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l315_1) begin
                  selectReadFifo_1 <= (selectReadFifo_1 + _zz_selectReadFifo_1_62);
                end
              end
            end
          end
          if(when_ArraySlice_l240_2) begin
            if(when_ArraySlice_l246_2) begin
              if(when_ArraySlice_l247_2) begin
                if(when_ArraySlice_l248_2) begin
                  selectReadFifo_2 <= (_zz_selectReadFifo_2_32 + _zz_selectReadFifo_2_34);
                end else begin
                  if(when_ArraySlice_l251_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + _zz_selectReadFifo_2_36);
                  end
                end
              end
              if(when_ArraySlice_l256_2) begin
                if(when_ArraySlice_l257_2) begin
                  if(when_ArraySlice_l259_2) begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_38 + _zz_selectReadFifo_2_40);
                  end else begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_42 + _zz_selectReadFifo_2_44);
                    if(when_ArraySlice_l265_2) begin
                      holdReadOp_2 <= 1'b1;
                    end
                    if(when_ArraySlice_l268_2) begin
                      allowPadding_2 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l272_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + _zz_selectReadFifo_2_46);
                  end
                end
              end
              if(when_ArraySlice_l276_2) begin
                if(when_ArraySlice_l277_2) begin
                  if(when_ArraySlice_l279_2) begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_48 + _zz_selectReadFifo_2_50);
                  end else begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_52 + _zz_selectReadFifo_2_54);
                    if(when_ArraySlice_l285_2) begin
                      holdReadOp_2 <= 1'b1;
                    end
                    if(when_ArraySlice_l288_2) begin
                      allowPadding_2 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l292_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + _zz_selectReadFifo_2_56);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l301_2) begin
              if(when_ArraySlice_l303_2) begin
                if(when_ArraySlice_l304_2) begin
                  selectReadFifo_2 <= (_zz_selectReadFifo_2_58 + _zz_selectReadFifo_2_60);
                end else begin
                  selectReadFifo_2 <= 6'h0;
                  readAround_2 <= (! readAround_2);
                  if(when_ArraySlice_l311_2) begin
                    holdReadOp_2 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l315_2) begin
                  selectReadFifo_2 <= (selectReadFifo_2 + _zz_selectReadFifo_2_62);
                end
              end
            end
          end
          if(when_ArraySlice_l240_3) begin
            if(when_ArraySlice_l246_3) begin
              if(when_ArraySlice_l247_3) begin
                if(when_ArraySlice_l248_3) begin
                  selectReadFifo_3 <= (_zz_selectReadFifo_3_32 + _zz_selectReadFifo_3_34);
                end else begin
                  if(when_ArraySlice_l251_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + _zz_selectReadFifo_3_36);
                  end
                end
              end
              if(when_ArraySlice_l256_3) begin
                if(when_ArraySlice_l257_3) begin
                  if(when_ArraySlice_l259_3) begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_38 + _zz_selectReadFifo_3_40);
                  end else begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_42 + _zz_selectReadFifo_3_44);
                    if(when_ArraySlice_l265_3) begin
                      holdReadOp_3 <= 1'b1;
                    end
                    if(when_ArraySlice_l268_3) begin
                      allowPadding_3 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l272_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + _zz_selectReadFifo_3_46);
                  end
                end
              end
              if(when_ArraySlice_l276_3) begin
                if(when_ArraySlice_l277_3) begin
                  if(when_ArraySlice_l279_3) begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_48 + _zz_selectReadFifo_3_50);
                  end else begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_52 + _zz_selectReadFifo_3_54);
                    if(when_ArraySlice_l285_3) begin
                      holdReadOp_3 <= 1'b1;
                    end
                    if(when_ArraySlice_l288_3) begin
                      allowPadding_3 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l292_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + _zz_selectReadFifo_3_56);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l301_3) begin
              if(when_ArraySlice_l303_3) begin
                if(when_ArraySlice_l304_3) begin
                  selectReadFifo_3 <= (_zz_selectReadFifo_3_58 + _zz_selectReadFifo_3_60);
                end else begin
                  selectReadFifo_3 <= 6'h0;
                  readAround_3 <= (! readAround_3);
                  if(when_ArraySlice_l311_3) begin
                    holdReadOp_3 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l315_3) begin
                  selectReadFifo_3 <= (selectReadFifo_3 + _zz_selectReadFifo_3_62);
                end
              end
            end
          end
          if(when_ArraySlice_l240_4) begin
            if(when_ArraySlice_l246_4) begin
              if(when_ArraySlice_l247_4) begin
                if(when_ArraySlice_l248_4) begin
                  selectReadFifo_4 <= (_zz_selectReadFifo_4_32 + _zz_selectReadFifo_4_34);
                end else begin
                  if(when_ArraySlice_l251_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + _zz_selectReadFifo_4_36);
                  end
                end
              end
              if(when_ArraySlice_l256_4) begin
                if(when_ArraySlice_l257_4) begin
                  if(when_ArraySlice_l259_4) begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_38 + _zz_selectReadFifo_4_40);
                  end else begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_42 + _zz_selectReadFifo_4_44);
                    if(when_ArraySlice_l265_4) begin
                      holdReadOp_4 <= 1'b1;
                    end
                    if(when_ArraySlice_l268_4) begin
                      allowPadding_4 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l272_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + _zz_selectReadFifo_4_46);
                  end
                end
              end
              if(when_ArraySlice_l276_4) begin
                if(when_ArraySlice_l277_4) begin
                  if(when_ArraySlice_l279_4) begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_48 + _zz_selectReadFifo_4_50);
                  end else begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_52 + _zz_selectReadFifo_4_54);
                    if(when_ArraySlice_l285_4) begin
                      holdReadOp_4 <= 1'b1;
                    end
                    if(when_ArraySlice_l288_4) begin
                      allowPadding_4 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l292_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + _zz_selectReadFifo_4_56);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l301_4) begin
              if(when_ArraySlice_l303_4) begin
                if(when_ArraySlice_l304_4) begin
                  selectReadFifo_4 <= (_zz_selectReadFifo_4_58 + _zz_selectReadFifo_4_60);
                end else begin
                  selectReadFifo_4 <= 6'h0;
                  readAround_4 <= (! readAround_4);
                  if(when_ArraySlice_l311_4) begin
                    holdReadOp_4 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l315_4) begin
                  selectReadFifo_4 <= (selectReadFifo_4 + _zz_selectReadFifo_4_62);
                end
              end
            end
          end
          if(when_ArraySlice_l240_5) begin
            if(when_ArraySlice_l246_5) begin
              if(when_ArraySlice_l247_5) begin
                if(when_ArraySlice_l248_5) begin
                  selectReadFifo_5 <= (_zz_selectReadFifo_5_32 + _zz_selectReadFifo_5_34);
                end else begin
                  if(when_ArraySlice_l251_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + _zz_selectReadFifo_5_36);
                  end
                end
              end
              if(when_ArraySlice_l256_5) begin
                if(when_ArraySlice_l257_5) begin
                  if(when_ArraySlice_l259_5) begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_38 + _zz_selectReadFifo_5_40);
                  end else begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_42 + _zz_selectReadFifo_5_44);
                    if(when_ArraySlice_l265_5) begin
                      holdReadOp_5 <= 1'b1;
                    end
                    if(when_ArraySlice_l268_5) begin
                      allowPadding_5 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l272_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + _zz_selectReadFifo_5_46);
                  end
                end
              end
              if(when_ArraySlice_l276_5) begin
                if(when_ArraySlice_l277_5) begin
                  if(when_ArraySlice_l279_5) begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_48 + _zz_selectReadFifo_5_50);
                  end else begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_52 + _zz_selectReadFifo_5_54);
                    if(when_ArraySlice_l285_5) begin
                      holdReadOp_5 <= 1'b1;
                    end
                    if(when_ArraySlice_l288_5) begin
                      allowPadding_5 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l292_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + _zz_selectReadFifo_5_56);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l301_5) begin
              if(when_ArraySlice_l303_5) begin
                if(when_ArraySlice_l304_5) begin
                  selectReadFifo_5 <= (_zz_selectReadFifo_5_58 + _zz_selectReadFifo_5_60);
                end else begin
                  selectReadFifo_5 <= 6'h0;
                  readAround_5 <= (! readAround_5);
                  if(when_ArraySlice_l311_5) begin
                    holdReadOp_5 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l315_5) begin
                  selectReadFifo_5 <= (selectReadFifo_5 + _zz_selectReadFifo_5_62);
                end
              end
            end
          end
          if(when_ArraySlice_l240_6) begin
            if(when_ArraySlice_l246_6) begin
              if(when_ArraySlice_l247_6) begin
                if(when_ArraySlice_l248_6) begin
                  selectReadFifo_6 <= (_zz_selectReadFifo_6_32 + _zz_selectReadFifo_6_34);
                end else begin
                  if(when_ArraySlice_l251_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + _zz_selectReadFifo_6_36);
                  end
                end
              end
              if(when_ArraySlice_l256_6) begin
                if(when_ArraySlice_l257_6) begin
                  if(when_ArraySlice_l259_6) begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_38 + _zz_selectReadFifo_6_40);
                  end else begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_42 + _zz_selectReadFifo_6_44);
                    if(when_ArraySlice_l265_6) begin
                      holdReadOp_6 <= 1'b1;
                    end
                    if(when_ArraySlice_l268_6) begin
                      allowPadding_6 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l272_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + _zz_selectReadFifo_6_46);
                  end
                end
              end
              if(when_ArraySlice_l276_6) begin
                if(when_ArraySlice_l277_6) begin
                  if(when_ArraySlice_l279_6) begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_48 + _zz_selectReadFifo_6_50);
                  end else begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_52 + _zz_selectReadFifo_6_54);
                    if(when_ArraySlice_l285_6) begin
                      holdReadOp_6 <= 1'b1;
                    end
                    if(when_ArraySlice_l288_6) begin
                      allowPadding_6 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l292_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + _zz_selectReadFifo_6_56);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l301_6) begin
              if(when_ArraySlice_l303_6) begin
                if(when_ArraySlice_l304_6) begin
                  selectReadFifo_6 <= (_zz_selectReadFifo_6_58 + _zz_selectReadFifo_6_60);
                end else begin
                  selectReadFifo_6 <= 6'h0;
                  readAround_6 <= (! readAround_6);
                  if(when_ArraySlice_l311_6) begin
                    holdReadOp_6 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l315_6) begin
                  selectReadFifo_6 <= (selectReadFifo_6 + _zz_selectReadFifo_6_62);
                end
              end
            end
          end
          if(when_ArraySlice_l240_7) begin
            if(when_ArraySlice_l246_7) begin
              if(when_ArraySlice_l247_7) begin
                if(when_ArraySlice_l248_7) begin
                  selectReadFifo_7 <= (_zz_selectReadFifo_7_32 + _zz_selectReadFifo_7_34);
                end else begin
                  if(when_ArraySlice_l251_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + _zz_selectReadFifo_7_36);
                  end
                end
              end
              if(when_ArraySlice_l256_7) begin
                if(when_ArraySlice_l257_7) begin
                  if(when_ArraySlice_l259_7) begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_38 + _zz_selectReadFifo_7_40);
                  end else begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_42 + _zz_selectReadFifo_7_44);
                    if(when_ArraySlice_l265_7) begin
                      holdReadOp_7 <= 1'b1;
                    end
                    if(when_ArraySlice_l268_7) begin
                      allowPadding_7 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l272_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + _zz_selectReadFifo_7_46);
                  end
                end
              end
              if(when_ArraySlice_l276_7) begin
                if(when_ArraySlice_l277_7) begin
                  if(when_ArraySlice_l279_7) begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_48 + _zz_selectReadFifo_7_50);
                  end else begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_52 + _zz_selectReadFifo_7_54);
                    if(when_ArraySlice_l285_7) begin
                      holdReadOp_7 <= 1'b1;
                    end
                    if(when_ArraySlice_l288_7) begin
                      allowPadding_7 <= 1'b0;
                    end
                  end
                end else begin
                  if(when_ArraySlice_l292_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + _zz_selectReadFifo_7_56);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l301_7) begin
              if(when_ArraySlice_l303_7) begin
                if(when_ArraySlice_l304_7) begin
                  selectReadFifo_7 <= (_zz_selectReadFifo_7_58 + _zz_selectReadFifo_7_60);
                end else begin
                  selectReadFifo_7 <= 6'h0;
                  readAround_7 <= (! readAround_7);
                  if(when_ArraySlice_l311_7) begin
                    holdReadOp_7 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l315_7) begin
                  selectReadFifo_7 <= (selectReadFifo_7 + _zz_selectReadFifo_7_62);
                end
              end
            end
          end
          if(when_ArraySlice_l333) begin
            if(when_ArraySlice_l338) begin
              if(when_ArraySlice_l339) begin
                selectWriteFifo <= 6'h0;
                writeAround <= (! writeAround);
              end else begin
                selectWriteFifo <= (selectWriteFifo + _zz_selectWriteFifo_2);
              end
            end
          end
          if(when_ArraySlice_l350) begin
            holdReadOp_0 <= 1'b0;
            holdReadOp_1 <= 1'b0;
            holdReadOp_2 <= 1'b0;
            holdReadOp_3 <= 1'b0;
            holdReadOp_4 <= 1'b0;
            holdReadOp_5 <= 1'b0;
            holdReadOp_6 <= 1'b0;
            holdReadOp_7 <= 1'b0;
          end
          if(when_ArraySlice_l358) begin
            if(when_ArraySlice_l361) begin
              allowPadding_0 <= 1'b1;
            end
            if(when_ArraySlice_l361_1) begin
              allowPadding_1 <= 1'b1;
            end
            if(when_ArraySlice_l361_2) begin
              allowPadding_2 <= 1'b1;
            end
            if(when_ArraySlice_l361_3) begin
              allowPadding_3 <= 1'b1;
            end
            if(when_ArraySlice_l361_4) begin
              allowPadding_4 <= 1'b1;
            end
            if(when_ArraySlice_l361_5) begin
              allowPadding_5 <= 1'b1;
            end
            if(when_ArraySlice_l361_6) begin
              allowPadding_6 <= 1'b1;
            end
            if(when_ArraySlice_l361_7) begin
              allowPadding_7 <= 1'b1;
            end
          end
        end
        default : begin
        end
      endcase
    end
  end


endmodule

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

module StreamFifo (
  input               io_push_valid,
  output              io_push_ready,
  input      [31:0]   io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [31:0]   io_pop_payload,
  input               io_flush,
  output     [6:0]    io_occupancy,
  output     [6:0]    io_availability,
  input               clk,
  input               resetn
);

  reg        [31:0]   _zz_logic_ram_port0;
  wire       [5:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [5:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [5:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [5:0]    logic_pushPtr_valueNext;
  reg        [5:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [5:0]    logic_popPtr_valueNext;
  reg        [5:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l946;
  wire       [5:0]    logic_ptrDif;
  reg [31:0] logic_ram [0:63];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {5'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {5'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= io_push_payload;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 6'h3f);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 6'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 6'h3f);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 6'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l946 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      logic_pushPtr_value <= 6'h0;
      logic_popPtr_value <= 6'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l946) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule
